module priority_mux(
    \p[0] ,
    \p[1] ,
    \p[2] ,
    \p[3] ,
    \p[4] ,
    \p[5] ,
    \p[6] ,
    \p[7] ,
    \p[8] ,
    \p[9] ,
    \p[10] ,
    \p[11] ,
    \p[12] ,
    \p[13] ,
    \p[14] ,
    \p[15] ,
    \p[16] ,
    \p[17] ,
    \p[18] ,
    \p[19] ,
    \p[20] ,
    \p[21] ,
    \p[22] ,
    \p[23] ,
    \p[24] ,
    \p[25] ,
    \p[26] ,
    \p[27] ,
    \p[28] ,
    \p[29] ,
    \p[30] ,
    \p[31] ,
    \p[32] ,
    \p[33] ,
    \p[34] ,
    \p[35] ,
    \p[36] ,
    \p[37] ,
    \p[38] ,
    \p[39] ,
    \p[40] ,
    \p[41] ,
    \p[42] ,
    \p[43] ,
    \p[44] ,
    \p[45] ,
    \p[46] ,
    \p[47] ,
    \p[48] ,
    \p[49] ,
    \p[50] ,
    \p[51] ,
    \p[52] ,
    \p[53] ,
    \p[54] ,
    \p[55] ,
    \p[56] ,
    \p[57] ,
    \p[58] ,
    \p[59] ,
    \p[60] ,
    \p[61] ,
    \p[62] ,
    \p[63] ,
    \p[64] ,
    \p[65] ,
    \p[66] ,
    \p[67] ,
    \p[68] ,
    \p[69] ,
    \p[70] ,
    \p[71] ,
    \p[72] ,
    \p[73] ,
    \p[74] ,
    \p[75] ,
    \p[76] ,
    \p[77] ,
    \p[78] ,
    \p[79] ,
    \p[80] ,
    \p[81] ,
    \p[82] ,
    \p[83] ,
    \p[84] ,
    \p[85] ,
    \p[86] ,
    \p[87] ,
    \p[88] ,
    \p[89] ,
    \p[90] ,
    \p[91] ,
    \p[92] ,
    \p[93] ,
    \p[94] ,
    \p[95] ,
    \p[96] ,
    \p[97] ,
    \p[98] ,
    \p[99] ,
    \p[100] ,
    \p[101] ,
    \p[102] ,
    \p[103] ,
    \p[104] ,
    \p[105] ,
    \p[106] ,
    \p[107] ,
    \p[108] ,
    \p[109] ,
    \p[110] ,
    \p[111] ,
    \p[112] ,
    \p[113] ,
    \p[114] ,
    \p[115] ,
    \p[116] ,
    \p[117] ,
    \p[118] ,
    \p[119] ,
    \p[120] ,
    \p[121] ,
    \p[122] ,
    \p[123] ,
    \p[124] ,
    \p[125] ,
    \p[126] ,
    \p[127] ,
    \p[128] ,
    \p[129] ,
    \p[130] ,
    \p[131] ,
    \p[132] ,
    \p[133] ,
    \p[134] ,
    \p[135] ,
    \p[136] ,
    \p[137] ,
    \p[138] ,
    \p[139] ,
    \p[140] ,
    \p[141] ,
    \p[142] ,
    \p[143] ,
    \p[144] ,
    \p[145] ,
    \p[146] ,
    \p[147] ,
    \p[148] ,
    \p[149] ,
    \p[150] ,
    \p[151] ,
    \p[152] ,
    \p[153] ,
    \p[154] ,
    \p[155] ,
    \p[156] ,
    \p[157] ,
    \p[158] ,
    \p[159] ,
    \p[160] ,
    \p[161] ,
    \p[162] ,
    \p[163] ,
    \p[164] ,
    \p[165] ,
    \p[166] ,
    \p[167] ,
    \p[168] ,
    \p[169] ,
    \p[170] ,
    \p[171] ,
    \p[172] ,
    \p[173] ,
    \p[174] ,
    \p[175] ,
    \p[176] ,
    \p[177] ,
    \p[178] ,
    \p[179] ,
    \p[180] ,
    \p[181] ,
    \p[182] ,
    \p[183] ,
    \p[184] ,
    \p[185] ,
    \p[186] ,
    \p[187] ,
    \p[188] ,
    \p[189] ,
    \p[190] ,
    \p[191] ,
    \p[192] ,
    \p[193] ,
    \p[194] ,
    \p[195] ,
    \p[196] ,
    \p[197] ,
    \p[198] ,
    \p[199] ,
    \p[200] ,
    \p[201] ,
    \p[202] ,
    \p[203] ,
    \p[204] ,
    \p[205] ,
    \p[206] ,
    \p[207] ,
    \p[208] ,
    \p[209] ,
    \p[210] ,
    \p[211] ,
    \p[212] ,
    \p[213] ,
    \p[214] ,
    \p[215] ,
    \p[216] ,
    \p[217] ,
    \p[218] ,
    \p[219] ,
    \p[220] ,
    \p[221] ,
    \p[222] ,
    \p[223] ,
    \p[224] ,
    \p[225] ,
    \p[226] ,
    \p[227] ,
    \p[228] ,
    \p[229] ,
    \p[230] ,
    \p[231] ,
    \p[232] ,
    \p[233] ,
    \p[234] ,
    \p[235] ,
    \p[236] ,
    \p[237] ,
    \p[238] ,
    \p[239] ,
    \p[240] ,
    \p[241] ,
    \p[242] ,
    \p[243] ,
    \p[244] ,
    \p[245] ,
    \p[246] ,
    \p[247] ,
    \p[248] ,
    \p[249] ,
    \p[250] ,
    \p[251] ,
    \p[252] ,
    \p[253] ,
    \p[254] ,
    \p[255] ,
    \v[0] ,
    \v[1] ,
    \v[2] ,
    \v[3] ,
    \v[4] ,
    \v[5] ,
    \v[6] ,
    \v[7] ,
    \v[8] ,
    \v[9] ,
    \v[10] ,
    \v[11] ,
    \v[12] ,
    \v[13] ,
    \v[14] ,
    \v[15] ,
    \v[16] ,
    \v[17] ,
    \v[18] ,
    \v[19] ,
    \v[20] ,
    \v[21] ,
    \v[22] ,
    \v[23] ,
    \v[24] ,
    \v[25] ,
    \v[26] ,
    \v[27] ,
    \v[28] ,
    \v[29] ,
    \v[30] ,
    \v[31] ,
    \v[32] ,
    \v[33] ,
    \v[34] ,
    \v[35] ,
    \v[36] ,
    \v[37] ,
    \v[38] ,
    \v[39] ,
    \v[40] ,
    \v[41] ,
    \v[42] ,
    \v[43] ,
    \v[44] ,
    \v[45] ,
    \v[46] ,
    \v[47] ,
    \v[48] ,
    \v[49] ,
    \v[50] ,
    \v[51] ,
    \v[52] ,
    \v[53] ,
    \v[54] ,
    \v[55] ,
    \v[56] ,
    \v[57] ,
    \v[58] ,
    \v[59] ,
    \v[60] ,
    \v[61] ,
    \v[62] ,
    \v[63] ,
    \v[64] ,
    \v[65] ,
    \v[66] ,
    \v[67] ,
    \v[68] ,
    \v[69] ,
    \v[70] ,
    \v[71] ,
    \v[72] ,
    \v[73] ,
    \v[74] ,
    \v[75] ,
    \v[76] ,
    \v[77] ,
    \v[78] ,
    \v[79] ,
    \v[80] ,
    \v[81] ,
    \v[82] ,
    \v[83] ,
    \v[84] ,
    \v[85] ,
    \v[86] ,
    \v[87] ,
    \v[88] ,
    \v[89] ,
    \v[90] ,
    \v[91] ,
    \v[92] ,
    \v[93] ,
    \v[94] ,
    \v[95] ,
    \v[96] ,
    \v[97] ,
    \v[98] ,
    \v[99] ,
    \v[100] ,
    \v[101] ,
    \v[102] ,
    \v[103] ,
    \v[104] ,
    \v[105] ,
    \v[106] ,
    \v[107] ,
    \v[108] ,
    \v[109] ,
    \v[110] ,
    \v[111] ,
    \v[112] ,
    \v[113] ,
    \v[114] ,
    \v[115] ,
    \v[116] ,
    \v[117] ,
    \v[118] ,
    \v[119] ,
    \v[120] ,
    \v[121] ,
    \v[122] ,
    \v[123] ,
    \v[124] ,
    \v[125] ,
    \v[126] ,
    \v[127] ,
    \v[128] ,
    \v[129] ,
    \v[130] ,
    \v[131] ,
    \v[132] ,
    \v[133] ,
    \v[134] ,
    \v[135] ,
    \v[136] ,
    \v[137] ,
    \v[138] ,
    \v[139] ,
    \v[140] ,
    \v[141] ,
    \v[142] ,
    \v[143] ,
    \v[144] ,
    \v[145] ,
    \v[146] ,
    \v[147] ,
    \v[148] ,
    \v[149] ,
    \v[150] ,
    \v[151] ,
    \v[152] ,
    \v[153] ,
    \v[154] ,
    \v[155] ,
    \v[156] ,
    \v[157] ,
    \v[158] ,
    \v[159] ,
    \v[160] ,
    \v[161] ,
    \v[162] ,
    \v[163] ,
    \v[164] ,
    \v[165] ,
    \v[166] ,
    \v[167] ,
    \v[168] ,
    \v[169] ,
    \v[170] ,
    \v[171] ,
    \v[172] ,
    \v[173] ,
    \v[174] ,
    \v[175] ,
    \v[176] ,
    \v[177] ,
    \v[178] ,
    \v[179] ,
    \v[180] ,
    \v[181] ,
    \v[182] ,
    \v[183] ,
    \v[184] ,
    \v[185] ,
    \v[186] ,
    \v[187] ,
    \v[188] ,
    \v[189] ,
    \v[190] ,
    \v[191] ,
    \v[192] ,
    \v[193] ,
    \v[194] ,
    \v[195] ,
    \v[196] ,
    \v[197] ,
    \v[198] ,
    \v[199] ,
    \v[200] ,
    \v[201] ,
    \v[202] ,
    \v[203] ,
    \v[204] ,
    \v[205] ,
    \v[206] ,
    \v[207] ,
    \v[208] ,
    \v[209] ,
    \v[210] ,
    \v[211] ,
    \v[212] ,
    \v[213] ,
    \v[214] ,
    \v[215] ,
    \v[216] ,
    \v[217] ,
    \v[218] ,
    \v[219] ,
    \v[220] ,
    \v[221] ,
    \v[222] ,
    \v[223] ,
    \v[224] ,
    \v[225] ,
    \v[226] ,
    \v[227] ,
    \v[228] ,
    \v[229] ,
    \v[230] ,
    \v[231] ,
    \v[232] ,
    \v[233] ,
    \v[234] ,
    \v[235] ,
    \v[236] ,
    \v[237] ,
    \v[238] ,
    \v[239] ,
    \v[240] ,
    \v[241] ,
    \v[242] ,
    \v[243] ,
    \v[244] ,
    \v[245] ,
    \v[246] ,
    \v[247] ,
    \v[248] ,
    \v[249] ,
    \v[250] ,
    \v[251] ,
    \v[252] ,
    \v[253] ,
    \v[254] ,
    \v[255] ,
    pp,
    vv,
    clk
);
    input clk;
    input \p[0] ;
    input \p[1] ;
    input \p[2] ;
    input \p[3] ;
    input \p[4] ;
    input \p[5] ;
    input \p[6] ;
    input \p[7] ;
    input \p[8] ;
    input \p[9] ;
    input \p[10] ;
    input \p[11] ;
    input \p[12] ;
    input \p[13] ;
    input \p[14] ;
    input \p[15] ;
    input \p[16] ;
    input \p[17] ;
    input \p[18] ;
    input \p[19] ;
    input \p[20] ;
    input \p[21] ;
    input \p[22] ;
    input \p[23] ;
    input \p[24] ;
    input \p[25] ;
    input \p[26] ;
    input \p[27] ;
    input \p[28] ;
    input \p[29] ;
    input \p[30] ;
    input \p[31] ;
    input \p[32] ;
    input \p[33] ;
    input \p[34] ;
    input \p[35] ;
    input \p[36] ;
    input \p[37] ;
    input \p[38] ;
    input \p[39] ;
    input \p[40] ;
    input \p[41] ;
    input \p[42] ;
    input \p[43] ;
    input \p[44] ;
    input \p[45] ;
    input \p[46] ;
    input \p[47] ;
    input \p[48] ;
    input \p[49] ;
    input \p[50] ;
    input \p[51] ;
    input \p[52] ;
    input \p[53] ;
    input \p[54] ;
    input \p[55] ;
    input \p[56] ;
    input \p[57] ;
    input \p[58] ;
    input \p[59] ;
    input \p[60] ;
    input \p[61] ;
    input \p[62] ;
    input \p[63] ;
    input \p[64] ;
    input \p[65] ;
    input \p[66] ;
    input \p[67] ;
    input \p[68] ;
    input \p[69] ;
    input \p[70] ;
    input \p[71] ;
    input \p[72] ;
    input \p[73] ;
    input \p[74] ;
    input \p[75] ;
    input \p[76] ;
    input \p[77] ;
    input \p[78] ;
    input \p[79] ;
    input \p[80] ;
    input \p[81] ;
    input \p[82] ;
    input \p[83] ;
    input \p[84] ;
    input \p[85] ;
    input \p[86] ;
    input \p[87] ;
    input \p[88] ;
    input \p[89] ;
    input \p[90] ;
    input \p[91] ;
    input \p[92] ;
    input \p[93] ;
    input \p[94] ;
    input \p[95] ;
    input \p[96] ;
    input \p[97] ;
    input \p[98] ;
    input \p[99] ;
    input \p[100] ;
    input \p[101] ;
    input \p[102] ;
    input \p[103] ;
    input \p[104] ;
    input \p[105] ;
    input \p[106] ;
    input \p[107] ;
    input \p[108] ;
    input \p[109] ;
    input \p[110] ;
    input \p[111] ;
    input \p[112] ;
    input \p[113] ;
    input \p[114] ;
    input \p[115] ;
    input \p[116] ;
    input \p[117] ;
    input \p[118] ;
    input \p[119] ;
    input \p[120] ;
    input \p[121] ;
    input \p[122] ;
    input \p[123] ;
    input \p[124] ;
    input \p[125] ;
    input \p[126] ;
    input \p[127] ;
    input \p[128] ;
    input \p[129] ;
    input \p[130] ;
    input \p[131] ;
    input \p[132] ;
    input \p[133] ;
    input \p[134] ;
    input \p[135] ;
    input \p[136] ;
    input \p[137] ;
    input \p[138] ;
    input \p[139] ;
    input \p[140] ;
    input \p[141] ;
    input \p[142] ;
    input \p[143] ;
    input \p[144] ;
    input \p[145] ;
    input \p[146] ;
    input \p[147] ;
    input \p[148] ;
    input \p[149] ;
    input \p[150] ;
    input \p[151] ;
    input \p[152] ;
    input \p[153] ;
    input \p[154] ;
    input \p[155] ;
    input \p[156] ;
    input \p[157] ;
    input \p[158] ;
    input \p[159] ;
    input \p[160] ;
    input \p[161] ;
    input \p[162] ;
    input \p[163] ;
    input \p[164] ;
    input \p[165] ;
    input \p[166] ;
    input \p[167] ;
    input \p[168] ;
    input \p[169] ;
    input \p[170] ;
    input \p[171] ;
    input \p[172] ;
    input \p[173] ;
    input \p[174] ;
    input \p[175] ;
    input \p[176] ;
    input \p[177] ;
    input \p[178] ;
    input \p[179] ;
    input \p[180] ;
    input \p[181] ;
    input \p[182] ;
    input \p[183] ;
    input \p[184] ;
    input \p[185] ;
    input \p[186] ;
    input \p[187] ;
    input \p[188] ;
    input \p[189] ;
    input \p[190] ;
    input \p[191] ;
    input \p[192] ;
    input \p[193] ;
    input \p[194] ;
    input \p[195] ;
    input \p[196] ;
    input \p[197] ;
    input \p[198] ;
    input \p[199] ;
    input \p[200] ;
    input \p[201] ;
    input \p[202] ;
    input \p[203] ;
    input \p[204] ;
    input \p[205] ;
    input \p[206] ;
    input \p[207] ;
    input \p[208] ;
    input \p[209] ;
    input \p[210] ;
    input \p[211] ;
    input \p[212] ;
    input \p[213] ;
    input \p[214] ;
    input \p[215] ;
    input \p[216] ;
    input \p[217] ;
    input \p[218] ;
    input \p[219] ;
    input \p[220] ;
    input \p[221] ;
    input \p[222] ;
    input \p[223] ;
    input \p[224] ;
    input \p[225] ;
    input \p[226] ;
    input \p[227] ;
    input \p[228] ;
    input \p[229] ;
    input \p[230] ;
    input \p[231] ;
    input \p[232] ;
    input \p[233] ;
    input \p[234] ;
    input \p[235] ;
    input \p[236] ;
    input \p[237] ;
    input \p[238] ;
    input \p[239] ;
    input \p[240] ;
    input \p[241] ;
    input \p[242] ;
    input \p[243] ;
    input \p[244] ;
    input \p[245] ;
    input \p[246] ;
    input \p[247] ;
    input \p[248] ;
    input \p[249] ;
    input \p[250] ;
    input \p[251] ;
    input \p[252] ;
    input \p[253] ;
    input \p[254] ;
    input \p[255] ;
    input \v[0] ;
    input \v[1] ;
    input \v[2] ;
    input \v[3] ;
    input \v[4] ;
    input \v[5] ;
    input \v[6] ;
    input \v[7] ;
    input \v[8] ;
    input \v[9] ;
    input \v[10] ;
    input \v[11] ;
    input \v[12] ;
    input \v[13] ;
    input \v[14] ;
    input \v[15] ;
    input \v[16] ;
    input \v[17] ;
    input \v[18] ;
    input \v[19] ;
    input \v[20] ;
    input \v[21] ;
    input \v[22] ;
    input \v[23] ;
    input \v[24] ;
    input \v[25] ;
    input \v[26] ;
    input \v[27] ;
    input \v[28] ;
    input \v[29] ;
    input \v[30] ;
    input \v[31] ;
    input \v[32] ;
    input \v[33] ;
    input \v[34] ;
    input \v[35] ;
    input \v[36] ;
    input \v[37] ;
    input \v[38] ;
    input \v[39] ;
    input \v[40] ;
    input \v[41] ;
    input \v[42] ;
    input \v[43] ;
    input \v[44] ;
    input \v[45] ;
    input \v[46] ;
    input \v[47] ;
    input \v[48] ;
    input \v[49] ;
    input \v[50] ;
    input \v[51] ;
    input \v[52] ;
    input \v[53] ;
    input \v[54] ;
    input \v[55] ;
    input \v[56] ;
    input \v[57] ;
    input \v[58] ;
    input \v[59] ;
    input \v[60] ;
    input \v[61] ;
    input \v[62] ;
    input \v[63] ;
    input \v[64] ;
    input \v[65] ;
    input \v[66] ;
    input \v[67] ;
    input \v[68] ;
    input \v[69] ;
    input \v[70] ;
    input \v[71] ;
    input \v[72] ;
    input \v[73] ;
    input \v[74] ;
    input \v[75] ;
    input \v[76] ;
    input \v[77] ;
    input \v[78] ;
    input \v[79] ;
    input \v[80] ;
    input \v[81] ;
    input \v[82] ;
    input \v[83] ;
    input \v[84] ;
    input \v[85] ;
    input \v[86] ;
    input \v[87] ;
    input \v[88] ;
    input \v[89] ;
    input \v[90] ;
    input \v[91] ;
    input \v[92] ;
    input \v[93] ;
    input \v[94] ;
    input \v[95] ;
    input \v[96] ;
    input \v[97] ;
    input \v[98] ;
    input \v[99] ;
    input \v[100] ;
    input \v[101] ;
    input \v[102] ;
    input \v[103] ;
    input \v[104] ;
    input \v[105] ;
    input \v[106] ;
    input \v[107] ;
    input \v[108] ;
    input \v[109] ;
    input \v[110] ;
    input \v[111] ;
    input \v[112] ;
    input \v[113] ;
    input \v[114] ;
    input \v[115] ;
    input \v[116] ;
    input \v[117] ;
    input \v[118] ;
    input \v[119] ;
    input \v[120] ;
    input \v[121] ;
    input \v[122] ;
    input \v[123] ;
    input \v[124] ;
    input \v[125] ;
    input \v[126] ;
    input \v[127] ;
    input \v[128] ;
    input \v[129] ;
    input \v[130] ;
    input \v[131] ;
    input \v[132] ;
    input \v[133] ;
    input \v[134] ;
    input \v[135] ;
    input \v[136] ;
    input \v[137] ;
    input \v[138] ;
    input \v[139] ;
    input \v[140] ;
    input \v[141] ;
    input \v[142] ;
    input \v[143] ;
    input \v[144] ;
    input \v[145] ;
    input \v[146] ;
    input \v[147] ;
    input \v[148] ;
    input \v[149] ;
    input \v[150] ;
    input \v[151] ;
    input \v[152] ;
    input \v[153] ;
    input \v[154] ;
    input \v[155] ;
    input \v[156] ;
    input \v[157] ;
    input \v[158] ;
    input \v[159] ;
    input \v[160] ;
    input \v[161] ;
    input \v[162] ;
    input \v[163] ;
    input \v[164] ;
    input \v[165] ;
    input \v[166] ;
    input \v[167] ;
    input \v[168] ;
    input \v[169] ;
    input \v[170] ;
    input \v[171] ;
    input \v[172] ;
    input \v[173] ;
    input \v[174] ;
    input \v[175] ;
    input \v[176] ;
    input \v[177] ;
    input \v[178] ;
    input \v[179] ;
    input \v[180] ;
    input \v[181] ;
    input \v[182] ;
    input \v[183] ;
    input \v[184] ;
    input \v[185] ;
    input \v[186] ;
    input \v[187] ;
    input \v[188] ;
    input \v[189] ;
    input \v[190] ;
    input \v[191] ;
    input \v[192] ;
    input \v[193] ;
    input \v[194] ;
    input \v[195] ;
    input \v[196] ;
    input \v[197] ;
    input \v[198] ;
    input \v[199] ;
    input \v[200] ;
    input \v[201] ;
    input \v[202] ;
    input \v[203] ;
    input \v[204] ;
    input \v[205] ;
    input \v[206] ;
    input \v[207] ;
    input \v[208] ;
    input \v[209] ;
    input \v[210] ;
    input \v[211] ;
    input \v[212] ;
    input \v[213] ;
    input \v[214] ;
    input \v[215] ;
    input \v[216] ;
    input \v[217] ;
    input \v[218] ;
    input \v[219] ;
    input \v[220] ;
    input \v[221] ;
    input \v[222] ;
    input \v[223] ;
    input \v[224] ;
    input \v[225] ;
    input \v[226] ;
    input \v[227] ;
    input \v[228] ;
    input \v[229] ;
    input \v[230] ;
    input \v[231] ;
    input \v[232] ;
    input \v[233] ;
    input \v[234] ;
    input \v[235] ;
    input \v[236] ;
    input \v[237] ;
    input \v[238] ;
    input \v[239] ;
    input \v[240] ;
    input \v[241] ;
    input \v[242] ;
    input \v[243] ;
    input \v[244] ;
    input \v[245] ;
    input \v[246] ;
    input \v[247] ;
    input \v[248] ;
    input \v[249] ;
    input \v[250] ;
    input \v[251] ;
    input \v[252] ;
    input \v[253] ;
    input \v[254] ;
    input \v[255] ;
    output pp;
    reg pp;
    output vv;
    reg vv;
    wire pp_ns;
    wire vv_ns;
    wire _0;
    wire _1;
    wire _2;
    wire _3;
    wire _4;
    wire _5;
    wire _6;
    wire _7;
    wire _8;
    wire _9;
    wire _10;
    wire _11;
    wire _12;
    wire _13;
    wire _14;
    wire _15;
    wire _16;
    wire _17;
    wire _18;
    wire _19;
    wire _20;
    wire _21;
    wire _22;
    wire _23;
    wire _24;
    wire _25;
    wire _26;
    wire _27;
    wire _28;
    wire _29;
    wire _30;
    wire _31;
    wire _32;
    wire _33;
    wire _34;
    wire _35;
    wire _36;
    wire _37;
    wire _38;
    wire _39;
    wire _40;
    wire _41;
    wire _42;
    wire _43;
    wire _44;
    wire _45;
    wire _46;
    wire _47;
    wire _48;
    wire _49;
    wire _50;
    wire _51;
    wire _52;
    wire _53;
    wire _54;
    wire _55;
    wire _56;
    wire _57;
    wire _58;
    wire _59;
    wire _60;
    wire _61;
    wire _62;
    wire _63;
    wire _64;
    wire _65;
    wire _66;
    wire _67;
    wire _68;
    wire _69;
    wire _70;
    wire _71;
    wire _72;
    wire _73;
    wire _74;
    wire _75;
    wire _76;
    wire _77;
    wire _78;
    wire _79;
    wire _80;
    wire _81;
    wire _82;
    wire _83;
    wire _84;
    wire _85;
    wire _86;
    wire _87;
    wire _88;
    wire _89;
    wire _90;
    wire _91;
    wire _92;
    wire _93;
    wire _94;
    wire _95;
    wire _96;
    wire _97;
    wire _98;
    wire _99;
    wire _100;
    wire _101;
    wire _102;
    wire _103;
    wire _104;
    wire _105;
    wire _106;
    wire _107;
    wire _108;
    wire _109;
    wire _110;
    wire _111;
    wire _112;
    wire _113;
    wire _114;
    wire _115;
    wire _116;
    wire _117;
    wire _118;
    wire _119;
    wire _120;
    wire _121;
    wire _122;
    wire _123;
    wire _124;
    wire _125;
    wire _126;
    wire _127;
    wire _128;
    wire _129;
    wire _130;
    wire _131;
    wire _132;
    wire _133;
    wire _134;
    wire _135;
    wire _136;
    wire _137;
    wire _138;
    wire _139;
    wire _140;
    wire _141;
    wire _142;
    wire _143;
    wire _144;
    wire _145;
    wire _146;
    wire _147;
    wire _148;
    wire _149;
    wire _150;
    wire _151;
    wire _152;
    wire _153;
    wire _154;
    wire _155;
    wire _156;
    wire _157;
    wire _158;
    wire _159;
    wire _160;
    wire _161;
    wire _162;
    wire _163;
    wire _164;
    wire _165;
    wire _166;
    wire _167;
    wire _168;
    wire _169;
    wire _170;
    wire _171;
    wire _172;
    wire _173;
    wire _174;
    wire _175;
    wire _176;
    wire _177;
    wire _178;
    wire _179;
    wire _180;
    wire _181;
    wire _182;
    wire _183;
    wire _184;
    wire _185;
    wire _186;
    wire _187;
    wire _188;
    wire _189;
    wire _190;
    wire _191;
    wire _192;
    wire _193;
    wire _194;
    wire _195;
    wire _196;
    wire _197;
    wire _198;
    wire _199;
    wire _200;
    wire _201;
    wire _202;
    wire _203;
    wire _204;
    wire _205;
    wire _206;
    wire _207;
    wire _208;
    wire _209;
    wire _210;
    wire _211;
    wire _212;
    wire _213;
    wire _214;
    wire _215;
    wire _216;
    wire _217;
    wire _218;
    wire _219;
    wire _220;
    wire _221;
    wire _222;
    wire _223;
    wire _224;
    wire _225;
    wire _226;
    wire _227;
    wire _228;
    wire _229;
    wire _230;
    wire _231;
    wire _232;
    wire _233;
    wire _234;
    wire _235;
    wire _236;
    wire _237;
    wire _238;
    wire _239;
    wire _240;
    wire _241;
    wire _242;
    wire _243;
    wire _244;
    wire _245;
    wire _246;
    wire _247;
    wire _248;
    wire _249;
    wire _250;
    wire _251;
    wire _252;
    wire _253;
    wire _254;
    wire _255;
    wire _256;
    wire _257;
    wire _258;
    wire _259;
    wire _260;
    wire _261;
    wire _262;
    wire _263;
    wire _264;
    wire _265;
    wire _266;
    wire _267;
    wire _268;
    wire _269;
    wire _270;
    wire _271;
    wire _272;
    wire _273;
    wire _274;
    wire _275;
    wire _276;
    wire _277;
    wire _278;
    wire _279;
    wire _280;
    wire _281;
    wire _282;
    wire _283;
    wire _284;
    wire _285;
    wire _286;
    wire _287;
    wire _288;
    wire _289;
    wire _290;
    wire _291;
    wire _292;
    wire _293;
    wire _294;
    wire _295;
    wire _296;
    wire _297;
    wire _298;
    wire _299;
    wire _300;
    wire _301;
    wire _302;
    wire _303;
    wire _304;
    wire _305;
    wire _306;
    wire _307;
    wire _308;
    wire _309;
    wire _310;
    wire _311;
    wire _312;
    wire _313;
    wire _314;
    wire _315;
    wire _316;
    wire _317;
    wire _318;
    wire _319;
    wire _320;
    wire _321;
    wire _322;
    wire _323;
    wire _324;
    wire _325;
    wire _326;
    wire _327;
    wire _328;
    wire _329;
    wire _330;
    wire _331;
    wire _332;
    wire _333;
    wire _334;
    wire _335;
    wire _336;
    wire _337;
    wire _338;
    wire _339;
    wire _340;
    wire _341;
    wire _342;
    wire _343;
    wire _344;
    wire _345;
    wire _346;
    wire _347;
    wire _348;
    wire _349;
    wire _350;
    wire _351;
    wire _352;
    wire _353;
    wire _354;
    wire _355;
    wire _356;
    wire _357;
    wire _358;
    wire _359;
    wire _360;
    wire _361;
    wire _362;
    wire _363;
    wire _364;
    wire _365;
    wire _366;
    wire _367;
    wire _368;
    wire _369;
    wire _370;
    wire _371;
    wire _372;
    wire _373;
    wire _374;
    wire _375;
    wire _376;
    wire _377;
    wire _378;
    wire _379;
    wire _380;
    wire _381;
    wire _382;
    wire _383;
    wire _384;
    wire _385;
    wire _386;
    wire _387;
    wire _388;
    wire _389;
    wire _390;
    wire _391;
    wire _392;
    wire _393;
    wire _394;
    wire _395;
    wire _396;
    wire _397;
    wire _398;
    wire _399;
    wire _400;
    wire _401;
    wire _402;
    wire _403;
    wire _404;
    wire _405;
    wire _406;
    wire _407;
    wire _408;
    wire _409;
    wire _410;
    wire _411;
    wire _412;
    wire _413;
    wire _414;
    wire _415;
    wire _416;
    wire _417;
    wire _418;
    wire _419;
    wire _420;
    wire _421;
    wire _422;
    wire _423;
    wire _424;
    wire _425;
    wire _426;
    wire _427;
    wire _428;
    wire _429;
    wire _430;
    wire _431;
    wire _432;
    wire _433;
    wire _434;
    wire _435;
    wire _436;
    wire _437;
    wire _438;
    wire _439;
    wire _440;
    wire _441;
    wire _442;
    wire _443;
    wire _444;
    wire _445;
    wire _446;
    wire _447;
    wire _448;
    wire _449;
    wire _450;
    wire _451;
    wire _452;
    wire _453;
    wire _454;
    wire _455;
    wire _456;
    wire _457;
    wire _458;
    wire _459;
    wire _460;
    wire _461;
    wire _462;
    wire _463;
    wire _464;
    wire _465;
    wire _466;
    wire _467;
    wire _468;
    wire _469;
    wire _470;
    wire _471;
    wire _472;
    wire _473;
    wire _474;
    wire _475;
    wire _476;
    wire _477;
    wire _478;
    wire _479;
    wire _480;
    wire _481;
    wire _482;
    wire _483;
    wire _484;
    wire _485;
    wire _486;
    wire _487;
    wire _488;
    wire _489;
    wire _490;
    wire _491;
    wire _492;
    wire _493;
    wire _494;
    wire _495;
    wire _496;
    wire _497;
    wire _498;
    wire _499;
    wire _500;
    wire _501;
    wire _502;
    wire _503;
    wire _504;
    wire _505;
    wire _506;
    wire _507;
    wire _508;
    wire _509;
    wire _510;
    wire _511;
    wire _512;
    wire _513;
    wire _514;
    wire _515;
    wire _516;
    wire _517;
    wire _518;
    wire _519;
    wire _520;
    wire _521;
    wire _522;
    wire _523;
    wire _524;
    wire _525;
    wire _526;
    wire _527;
    wire _528;
    wire _529;
    wire _530;
    wire _531;
    wire _532;
    wire _533;
    wire _534;
    wire _535;
    wire _536;
    wire _537;
    wire _538;
    wire _539;
    wire _540;
    wire _541;
    wire _542;
    wire _543;
    wire _544;
    wire _545;
    wire _546;
    wire _547;
    wire _548;
    wire _549;
    wire _550;
    wire _551;
    wire _552;
    wire _553;
    wire _554;
    wire _555;
    wire _556;
    wire _557;
    wire _558;
    wire _559;
    wire _560;
    wire _561;
    wire _562;
    wire _563;
    wire _564;
    wire _565;
    wire _566;
    wire _567;
    wire _568;
    wire _569;
    wire _570;
    wire _571;
    wire _572;
    wire _573;
    wire _574;
    wire _575;
    wire _576;
    wire _577;
    wire _578;
    wire _579;
    wire _580;
    wire _581;
    wire _582;
    wire _583;
    wire _584;
    wire _585;
    wire _586;
    wire _587;
    wire _588;
    wire _589;
    wire _590;
    wire _591;
    wire _592;
    wire _593;
    wire _594;
    wire _595;
    wire _596;
    wire _597;
    wire _598;
    wire _599;
    wire _600;
    wire _601;
    wire _602;
    wire _603;
    wire _604;
    wire _605;
    wire _606;
    wire _607;
    wire _608;
    wire _609;
    wire _610;
    wire _611;
    wire _612;
    wire _613;
    wire _614;
    wire _615;
    wire _616;
    wire _617;
    wire _618;
    wire _619;
    wire _620;
    wire _621;
    wire _622;
    wire _623;
    wire _624;
    wire _625;
    wire _626;
    wire _627;
    wire _628;
    wire _629;
    wire _630;
    wire _631;
    wire _632;
    wire _633;
    wire _634;
    wire _635;
    wire _636;
    wire _637;
    wire _638;
    wire _639;
    wire _640;
    wire _641;
    wire _642;
    wire _643;
    wire _644;
    wire _645;
    wire _646;
    wire _647;
    wire _648;
    wire _649;
    wire _650;
    wire _651;
    wire _652;
    wire _653;
    wire _654;
    wire _655;
    wire _656;
    wire _657;
    wire _658;
    wire _659;
    wire _660;
    wire _661;
    wire _662;
    wire _663;
    wire _664;
    wire _665;
    wire _666;
    wire _667;
    wire _668;
    wire _669;
    wire _670;
    wire _671;
    wire _672;
    wire _673;
    wire _674;
    wire _675;
    wire _676;
    wire _677;
    wire _678;
    wire _679;
    wire _680;
    wire _681;
    wire _682;
    wire _683;
    wire _684;
    wire _685;
    wire _686;
    wire _687;
    wire _688;
    wire _689;
    wire _690;
    wire _691;
    wire _692;
    wire _693;
    wire _694;
    wire _695;
    wire _696;
    wire _697;
    wire _698;
    wire _699;
    wire _700;
    wire _701;
    wire _702;
    wire _703;
    wire _704;
    wire _705;
    wire _706;
    wire _707;
    wire _708;
    wire _709;
    wire _710;
    wire _711;
    wire _712;
    wire _713;
    wire _714;
    wire _715;
    wire _716;
    wire _717;
    wire _718;
    wire _719;
    wire _720;
    wire _721;
    wire _722;
    wire _723;
    wire _724;
    wire _725;
    wire _726;
    wire _727;
    wire _728;
    wire _729;
    wire _730;
    wire _731;
    wire _732;
    wire _733;
    wire _734;
    wire _735;
    wire _736;
    wire _737;
    wire _738;
    wire _739;
    wire _740;
    wire _741;
    wire _742;
    wire _743;
    wire _744;
    wire _745;
    wire _746;
    wire _747;
    wire _748;
    wire _749;
    wire _750;
    wire _751;
    wire _752;
    wire _753;
    wire _754;
    wire _755;
    wire _756;
    wire _757;
    wire _758;
    wire _759;
    wire _760;
    wire _761;
    wire _762;
    wire _763;
    wire _764;
    wire _765;
    wire _766;
    wire _767;
    wire _768;
    wire _769;
    wire _770;
    wire _771;
    wire _772;
    wire _773;
    wire _774;
    wire _775;
    wire _776;
    wire _777;
    wire _778;
    wire _779;
    wire _780;
    wire _781;
    wire _782;
    wire _783;
    wire _784;
    wire _785;
    wire _786;
    wire _787;
    wire _788;
    wire _789;
    wire _790;
    wire _791;
    wire _792;
    wire _793;
    wire _794;
    wire _795;
    wire _796;
    wire _797;
    wire _798;
    wire _799;
    wire _800;
    wire _801;
    wire _802;
    wire _803;
    wire _804;
    wire _805;
    wire _806;
    wire _807;
    wire _808;
    wire _809;
    wire _810;
    wire _811;
    wire _812;
    wire _813;
    wire _814;
    wire _815;
    wire _816;
    wire _817;
    wire _818;
    wire _819;
    wire _820;
    wire _821;
    wire _822;
    wire _823;
    wire _824;
    wire _825;
    wire _826;
    wire _827;
    wire _828;
    wire _829;
    wire _830;
    wire _831;
    wire _832;
    wire _833;
    wire _834;
    wire _835;
    wire _836;
    wire _837;
    wire _838;
    wire _839;
    wire _840;
    wire _841;
    wire _842;
    wire _843;
    wire _844;
    wire _845;
    wire _846;
    wire _847;
    wire _848;
    wire _849;
    wire _850;
    wire _851;
    wire _852;
    wire _853;
    wire _854;
    wire _855;
    wire _856;
    wire _857;
    wire _858;
    wire _859;
    wire _860;
    wire _861;
    wire _862;
    wire _863;
    wire _864;
    wire _865;
    wire _866;
    wire _867;
    wire _868;
    wire _869;
    wire _870;
    wire _871;
    wire _872;
    wire _873;
    wire _874;
    wire _875;
    wire _876;
    wire _877;
    wire _878;
    wire _879;
    wire _880;
    wire _881;
    wire _882;
    wire _883;
    wire _884;
    wire _885;
    wire _886;
    wire _887;
    wire _888;
    wire _889;
    wire _890;
    wire _891;
    wire _892;
    wire _893;
    wire _894;
    wire _895;
    wire _896;
    wire _897;
    wire _898;
    wire _899;
    wire _900;
    wire _901;
    wire _902;
    wire _903;
    wire _904;
    wire _905;
    wire _906;
    wire _907;
    wire _908;
    wire _909;
    wire _910;
    wire _911;
    wire _912;
    wire _913;
    wire _914;
    wire _915;
    wire _916;
    wire _917;
    wire _918;
    wire _919;
    wire _920;
    wire _921;
    wire _922;
    wire _923;
    wire _924;
    wire _925;
    wire _926;
    wire _927;
    wire _928;
    wire _929;
    wire _930;
    wire _931;
    wire _932;
    wire _933;
    wire _934;
    wire _935;
    wire _936;
    wire _937;
    wire _938;
    wire _939;
    wire _940;
    wire _941;
    wire _942;
    wire _943;
    wire _944;
    wire _945;
    wire _946;
    wire _947;
    wire _948;
    wire _949;
    wire _950;
    wire _951;
    wire _952;
    wire _953;
    wire _954;
    wire _955;
    wire _956;
    wire _957;
    wire _958;
    wire _959;
    wire _960;
    wire _961;
    wire _962;
    wire _963;
    wire _964;
    wire _965;
    wire _966;
    wire _967;
    wire _968;
    wire _969;
    wire _970;
    wire _971;
    wire _972;
    wire _973;
    wire _974;
    wire _975;
    wire _976;
    wire _977;
    wire _978;
    wire _979;
    wire _980;
    wire _981;
    wire _982;
    wire _983;
    wire _984;
    wire _985;
    wire _986;
    wire _987;
    wire _988;
    wire _989;
    wire _990;
    wire _991;
    wire _992;
    wire _993;
    wire _994;
    wire _995;
    wire _996;
    wire _997;
    wire _998;
    wire _999;
    wire _1000;
    wire _1001;
    wire _1002;
    wire _1003;
    wire _1004;
    wire _1005;
    wire _1006;
    wire _1007;
    wire _1008;
    wire _1009;
    wire _1010;
    wire _1011;
    wire _1012;
    wire _1013;
    wire _1014;
    wire _1015;
    wire _1016;
    wire _1017;
    wire _1018;
    wire _1019;
    wire _1020;
    wire _1021;
    wire _1022;
    wire _1023;
    wire _1024;
    wire _1025;
    wire _1026;
    wire _1027;
    wire _1028;
    wire _1029;
    wire _1030;
    wire _1031;
    wire _1032;
    wire _1033;
    wire _1034;
    wire _1035;
    wire _1036;
    wire _1037;
    wire _1038;
    wire _1039;
    wire _1040;
    wire _1041;
    wire _1042;
    wire _1043;
    wire _1044;
    wire _1045;
    wire _1046;
    wire _1047;
    wire _1048;
    wire _1049;
    wire _1050;
    wire _1051;
    wire _1052;
    wire _1053;
    wire _1054;
    wire _1055;
    wire _1056;
    wire _1057;
    wire _1058;
    wire _1059;
    wire _1060;
    wire _1061;
    wire _1062;
    wire _1063;
    wire _1064;
    wire _1065;
    wire _1066;
    wire _1067;
    wire _1068;
    wire _1069;
    wire _1070;
    wire _1071;
    wire _1072;
    wire _1073;
    wire _1074;
    wire _1075;
    wire _1076;
    wire _1077;
    wire _1078;
    wire _1079;
    wire _1080;
    wire _1081;
    wire _1082;
    wire _1083;
    wire _1084;
    wire _1085;
    wire _1086;
    wire _1087;
    wire _1088;
    wire _1089;
    wire _1090;
    wire _1091;
    wire _1092;
    wire _1093;
    wire _1094;
    wire _1095;
    wire _1096;
    wire _1097;
    wire _1098;
    wire _1099;
    wire _1100;
    wire _1101;
    wire _1102;
    wire _1103;
    wire _1104;
    wire _1105;
    wire _1106;
    wire _1107;
    wire _1108;
    wire _1109;
    wire _1110;
    wire _1111;
    wire _1112;
    wire _1113;
    wire _1114;
    wire _1115;
    wire _1116;
    wire _1117;
    wire _1118;
    wire _1119;
    wire _1120;
    wire _1121;
    wire _1122;
    wire _1123;
    wire _1124;
    wire _1125;
    wire _1126;
    wire _1127;
    wire _1128;
    wire _1129;
    wire _1130;
    wire _1131;
    wire _1132;
    wire _1133;
    wire _1134;
    wire _1135;
    wire _1136;
    wire _1137;
    wire _1138;
    wire _1139;
    wire _1140;
    wire _1141;
    wire _1142;
    wire _1143;
    wire _1144;
    wire _1145;
    wire _1146;
    wire _1147;
    wire _1148;
    wire _1149;
    wire _1150;
    wire _1151;
    wire _1152;
    wire _1153;
    wire _1154;
    wire _1155;
    wire _1156;
    wire _1157;
    wire _1158;
    wire _1159;
    wire _1160;
    wire _1161;
    wire _1162;
    wire _1163;
    wire _1164;
    wire _1165;
    wire _1166;
    wire _1167;
    wire _1168;
    wire _1169;
    wire _1170;
    wire _1171;
    wire _1172;
    wire _1173;
    wire _1174;
    wire _1175;
    wire _1176;
    wire _1177;
    wire _1178;
    wire _1179;
    wire _1180;
    wire _1181;
    wire _1182;
    wire _1183;
    wire _1184;
    wire _1185;
    wire _1186;
    wire _1187;
    wire _1188;
    wire _1189;
    wire _1190;
    wire _1191;
    wire _1192;
    wire _1193;
    wire _1194;
    wire _1195;
    wire _1196;
    wire _1197;
    wire _1198;
    wire _1199;
    wire _1200;
    wire _1201;
    wire _1202;
    wire _1203;
    wire _1204;
    wire _1205;
    wire _1206;
    wire _1207;
    wire _1208;
    wire _1209;
    wire _1210;
    wire _1211;
    wire _1212;
    wire _1213;
    wire _1214;
    wire _1215;
    wire _1216;
    wire _1217;
    wire _1218;
    wire _1219;
    wire _1220;
    wire _1221;
    wire _1222;
    wire _1223;
    wire _1224;
    wire _1225;
    wire _1226;
    wire _1227;
    wire _1228;
    wire _1229;
    wire _1230;
    wire _1231;
    wire _1232;
    wire _1233;
    wire _1234;
    wire _1235;
    wire _1236;
    wire _1237;
    wire _1238;
    wire _1239;
    wire _1240;
    wire _1241;
    wire _1242;
    wire _1243;
    wire _1244;
    wire _1245;
    wire _1246;
    wire _1247;
    wire _1248;
    wire _1249;
    wire _1250;
    wire _1251;
    wire _1252;
    wire _1253;
    wire _1254;
    wire _1255;
    wire _1256;
    wire _1257;
    wire _1258;
    wire _1259;
    wire _1260;
    wire _1261;
    wire _1262;
    wire _1263;
    wire _1264;
    wire _1265;
    wire _1266;
    wire _1267;
    wire _1268;
    wire _1269;
    wire _1270;
    wire _1271;
    wire _1272;
    wire _1273;
    wire _1274;
    wire _1275;
    wire _1276;
    wire _1277;
    wire _1278;
    wire _1279;
    wire _1280;
    wire _1281;
    wire _1282;
    wire _1283;
    wire _1284;
    wire _1285;
    wire _1286;
    wire _1287;
    wire _1288;
    wire _1289;
    wire _1290;
    wire _1291;
    wire _1292;
    wire _1293;
    wire _1294;
    wire _1295;
    wire _1296;
    wire _1297;
    wire _1298;
    wire _1299;
    wire _1300;
    wire _1301;
    wire _1302;
    wire _1303;
    wire _1304;
    wire _1305;
    wire _1306;
    wire _1307;
    wire _1308;
    wire _1309;
    wire _1310;
    wire _1311;
    wire _1312;
    wire _1313;
    wire _1314;
    wire _1315;
    wire _1316;
    wire _1317;
    wire _1318;
    wire _1319;
    wire _1320;
    wire _1321;
    wire _1322;
    wire _1323;
    wire _1324;
    wire _1325;
    wire _1326;
    wire _1327;
    wire _1328;
    wire _1329;
    wire _1330;
    wire _1331;
    wire _1332;
    wire _1333;
    wire _1334;
    wire _1335;
    wire _1336;
    wire _1337;
    wire _1338;
    wire _1339;
    wire _1340;
    wire _1341;
    wire _1342;
    wire _1343;
    wire _1344;
    wire _1345;
    wire _1346;
    wire _1347;
    wire _1348;
    wire _1349;
    wire _1350;
    wire _1351;
    wire _1352;
    wire _1353;
    wire _1354;
    wire _1355;
    wire _1356;
    wire _1357;
    wire _1358;
    wire _1359;
    wire _1360;
    wire _1361;
    wire _1362;
    wire _1363;
    wire _1364;
    wire _1365;
    wire _1366;
    wire _1367;
    wire _1368;
    wire _1369;
    wire _1370;
    wire _1371;
    wire _1372;
    wire _1373;
    wire _1374;
    wire _1375;
    wire _1376;
    wire _1377;
    wire _1378;
    wire _1379;
    wire _1380;
    wire _1381;
    wire _1382;
    wire _1383;
    wire _1384;
    wire _1385;
    wire _1386;
    wire _1387;
    wire _1388;
    wire _1389;
    wire _1390;
    wire _1391;
    wire _1392;
    wire _1393;
    wire _1394;
    wire _1395;
    wire _1396;
    wire _1397;
    wire _1398;
    wire _1399;
    wire _1400;
    wire _1401;
    wire _1402;
    wire _1403;
    wire _1404;
    wire _1405;
    wire _1406;
    wire _1407;
    wire _1408;
    wire _1409;
    wire _1410;
    wire _1411;
    wire _1412;
    wire _1413;
    wire _1414;
    wire _1415;
    wire _1416;
    wire _1417;
    wire _1418;
    wire _1419;
    wire _1420;
    wire _1421;
    wire _1422;
    wire _1423;
    wire _1424;
    wire _1425;
    wire _1426;
    wire _1427;
    wire _1428;
    wire _1429;
    wire _1430;
    wire _1431;
    wire _1432;
    wire _1433;
    wire _1434;
    wire _1435;
    wire _1436;
    wire _1437;
    wire _1438;
    wire _1439;
    wire _1440;
    wire _1441;
    wire _1442;
    wire _1443;
    wire _1444;
    wire _1445;
    wire _1446;
    wire _1447;
    wire _1448;
    wire _1449;
    wire _1450;
    wire _1451;
    wire _1452;
    wire _1453;
    wire _1454;
    wire _1455;
    wire _1456;
    wire _1457;
    wire _1458;
    wire _1459;
    wire _1460;
    wire _1461;
    wire _1462;
    wire _1463;
    wire _1464;
    wire _1465;
    wire _1466;
    wire _1467;
    wire _1468;
    wire _1469;
    wire _1470;
    wire _1471;
    wire _1472;
    wire _1473;
    wire _1474;
    wire _1475;
    wire _1476;
    wire _1477;
    wire _1478;
    wire _1479;
    wire _1480;
    wire _1481;
    wire _1482;
    wire _1483;
    wire _1484;
    wire _1485;
    wire _1486;
    wire _1487;
    wire _1488;
    wire _1489;
    wire _1490;
    wire _1491;
    wire _1492;
    wire _1493;
    wire _1494;
    wire _1495;
    wire _1496;
    wire _1497;
    wire _1498;
    wire _1499;
    wire _1500;
    wire _1501;
    wire _1502;
    wire _1503;
    wire _1504;
    wire _1505;
    wire _1506;
    wire _1507;
    wire _1508;
    wire _1509;
    wire _1510;
    wire _1511;
    wire _1512;
    wire _1513;
    wire _1514;
    wire _1515;
    wire _1516;
    wire _1517;
    wire _1518;
    wire _1519;
    wire _1520;
    wire _1521;
    wire _1522;
    wire _1523;
    wire _1524;
    wire _1525;
    wire _1526;
    wire _1527;
    wire _1528;
    wire _1529;
    wire _1530;
    wire _1531;
    wire _1532;
    wire _1533;
    wire _1534;
    wire _1535;
    wire _1536;
    wire _1537;
    wire _1538;
    wire _1539;
    wire _1540;
    wire _1541;
    wire _1542;
    wire _1543;
    wire _1544;
    wire _1545;
    wire _1546;
    wire _1547;
    wire _1548;
    wire _1549;
    wire _1550;
    wire _1551;
    wire _1552;
    wire _1553;
    wire _1554;
    wire _1555;
    wire _1556;
    wire _1557;
    wire _1558;
    wire _1559;
    wire _1560;
    wire _1561;
    wire _1562;
    wire _1563;
    wire _1564;
    wire _1565;
    wire _1566;
    wire _1567;
    wire _1568;
    wire _1569;
    wire _1570;
    wire _1571;
    wire _1572;
    wire _1573;
    wire _1574;
    wire _1575;
    wire _1576;
    wire _1577;
    wire _1578;
    wire _1579;
    wire _1580;
    wire _1581;
    wire _1582;
    wire _1583;
    wire _1584;
    wire _1585;
    wire _1586;
    wire _1587;
    wire _1588;
    wire _1589;
    wire _1590;
    wire _1591;
    wire _1592;
    wire _1593;
    wire _1594;
    wire _1595;
    wire _1596;
    wire _1597;
    wire _1598;
    wire _1599;
    wire _1600;
    wire _1601;
    wire _1602;
    wire _1603;
    wire _1604;
    wire _1605;
    wire _1606;
    wire _1607;
    wire _1608;
    wire _1609;
    wire _1610;
    wire _1611;
    wire _1612;
    wire _1613;
    wire _1614;
    wire _1615;
    wire _1616;
    wire _1617;
    wire _1618;
    wire _1619;
    wire _1620;
    wire _1621;
    wire _1622;
    wire _1623;
    wire _1624;
    wire _1625;
    wire _1626;
    wire _1627;
    wire _1628;
    wire _1629;
    wire _1630;
    wire _1631;
    wire _1632;
    wire _1633;
    wire _1634;
    wire _1635;
    wire _1636;
    wire _1637;
    wire _1638;
    wire _1639;
    wire _1640;
    wire _1641;
    wire _1642;
    wire _1643;
    wire _1644;
    wire _1645;
    wire _1646;
    wire _1647;
    wire _1648;
    wire _1649;
    wire _1650;
    wire _1651;
    wire _1652;
    wire _1653;
    wire _1654;
    wire _1655;
    wire _1656;
    wire _1657;
    wire _1658;
    wire _1659;
    wire _1660;
    wire _1661;
    wire _1662;
    wire _1663;
    wire _1664;
    wire _1665;
    wire _1666;
    wire _1667;
    wire _1668;
    wire _1669;
    wire _1670;
    wire _1671;
    wire _1672;
    wire _1673;
    wire _1674;
    wire _1675;
    wire _1676;
    wire _1677;
    wire _1678;
    wire _1679;
    wire _1680;
    wire _1681;
    wire _1682;
    wire _1683;
    wire _1684;
    wire _1685;
    wire _1686;
    wire _1687;
    wire _1688;
    wire _1689;
    wire _1690;
    wire _1691;
    wire _1692;
    wire _1693;
    wire _1694;
    wire _1695;
    wire _1696;
    wire _1697;
    wire _1698;
    wire _1699;
    wire _1700;
    wire _1701;
    wire _1702;
    wire _1703;
    wire _1704;
    wire _1705;
    wire _1706;
    wire _1707;
    wire _1708;
    wire _1709;
    wire _1710;
    wire _1711;
    wire _1712;
    wire _1713;
    wire _1714;
    wire _1715;
    wire _1716;
    wire _1717;
    wire _1718;
    wire _1719;
    wire _1720;
    wire _1721;
    wire _1722;
    wire _1723;
    wire _1724;
    wire _1725;
    wire _1726;
    wire _1727;
    wire _1728;
    wire _1729;
    wire _1730;
    wire _1731;
    wire _1732;
    wire _1733;
    wire _1734;
    wire _1735;
    wire _1736;
    wire _1737;
    wire _1738;
    wire _1739;
    wire _1740;
    wire _1741;
    wire _1742;
    wire _1743;
    wire _1744;
    wire _1745;
    wire _1746;
    wire _1747;
    wire _1748;
    wire _1749;
    wire _1750;
    wire _1751;
    wire _1752;
    wire _1753;
    wire _1754;
    wire _1755;
    wire _1756;
    wire _1757;
    wire _1758;
    wire _1759;
    wire _1760;
    wire _1761;
    wire _1762;
    wire _1763;
    wire _1764;
    wire _1765;
    wire _1766;
    wire _1767;
    wire _1768;
    wire _1769;
    wire _1770;
    wire _1771;
    wire _1772;
    wire _1773;
    wire _1774;
    wire _1775;
    wire _1776;
    wire _1777;
    wire _1778;
    wire _1779;
    wire _1780;
    wire _1781;
    wire _1782;
    wire _1783;
    wire _1784;
    wire _1785;
    wire _1786;
    assign _0 = \p[0] ;
    assign _1 = \p[1] ;
    assign _2 = \p[2] ;
    assign _3 = \p[3] ;
    assign _4 = \p[4] ;
    assign _5 = \p[5] ;
    assign _6 = \p[6] ;
    assign _7 = \p[7] ;
    assign _8 = \p[8] ;
    assign _9 = \p[9] ;
    assign _10 = \p[10] ;
    assign _11 = \p[11] ;
    assign _12 = \p[12] ;
    assign _13 = \p[13] ;
    assign _14 = \p[14] ;
    assign _15 = \p[15] ;
    assign _16 = \p[16] ;
    assign _17 = \p[17] ;
    assign _18 = \p[18] ;
    assign _19 = \p[19] ;
    assign _20 = \p[20] ;
    assign _21 = \p[21] ;
    assign _22 = \p[22] ;
    assign _23 = \p[23] ;
    assign _24 = \p[24] ;
    assign _25 = \p[25] ;
    assign _26 = \p[26] ;
    assign _27 = \p[27] ;
    assign _28 = \p[28] ;
    assign _29 = \p[29] ;
    assign _30 = \p[30] ;
    assign _31 = \p[31] ;
    assign _32 = \p[32] ;
    assign _33 = \p[33] ;
    assign _34 = \p[34] ;
    assign _35 = \p[35] ;
    assign _36 = \p[36] ;
    assign _37 = \p[37] ;
    assign _38 = \p[38] ;
    assign _39 = \p[39] ;
    assign _40 = \p[40] ;
    assign _41 = \p[41] ;
    assign _42 = \p[42] ;
    assign _43 = \p[43] ;
    assign _44 = \p[44] ;
    assign _45 = \p[45] ;
    assign _46 = \p[46] ;
    assign _47 = \p[47] ;
    assign _48 = \p[48] ;
    assign _49 = \p[49] ;
    assign _50 = \p[50] ;
    assign _51 = \p[51] ;
    assign _52 = \p[52] ;
    assign _53 = \p[53] ;
    assign _54 = \p[54] ;
    assign _55 = \p[55] ;
    assign _56 = \p[56] ;
    assign _57 = \p[57] ;
    assign _58 = \p[58] ;
    assign _59 = \p[59] ;
    assign _60 = \p[60] ;
    assign _61 = \p[61] ;
    assign _62 = \p[62] ;
    assign _63 = \p[63] ;
    assign _64 = \p[64] ;
    assign _65 = \p[65] ;
    assign _66 = \p[66] ;
    assign _67 = \p[67] ;
    assign _68 = \p[68] ;
    assign _69 = \p[69] ;
    assign _70 = \p[70] ;
    assign _71 = \p[71] ;
    assign _72 = \p[72] ;
    assign _73 = \p[73] ;
    assign _74 = \p[74] ;
    assign _75 = \p[75] ;
    assign _76 = \p[76] ;
    assign _77 = \p[77] ;
    assign _78 = \p[78] ;
    assign _79 = \p[79] ;
    assign _80 = \p[80] ;
    assign _81 = \p[81] ;
    assign _82 = \p[82] ;
    assign _83 = \p[83] ;
    assign _84 = \p[84] ;
    assign _85 = \p[85] ;
    assign _86 = \p[86] ;
    assign _87 = \p[87] ;
    assign _88 = \p[88] ;
    assign _89 = \p[89] ;
    assign _90 = \p[90] ;
    assign _91 = \p[91] ;
    assign _92 = \p[92] ;
    assign _93 = \p[93] ;
    assign _94 = \p[94] ;
    assign _95 = \p[95] ;
    assign _96 = \p[96] ;
    assign _97 = \p[97] ;
    assign _98 = \p[98] ;
    assign _99 = \p[99] ;
    assign _100 = \p[100] ;
    assign _101 = \p[101] ;
    assign _102 = \p[102] ;
    assign _103 = \p[103] ;
    assign _104 = \p[104] ;
    assign _105 = \p[105] ;
    assign _106 = \p[106] ;
    assign _107 = \p[107] ;
    assign _108 = \p[108] ;
    assign _109 = \p[109] ;
    assign _110 = \p[110] ;
    assign _111 = \p[111] ;
    assign _112 = \p[112] ;
    assign _113 = \p[113] ;
    assign _114 = \p[114] ;
    assign _115 = \p[115] ;
    assign _116 = \p[116] ;
    assign _117 = \p[117] ;
    assign _118 = \p[118] ;
    assign _119 = \p[119] ;
    assign _120 = \p[120] ;
    assign _121 = \p[121] ;
    assign _122 = \p[122] ;
    assign _123 = \p[123] ;
    assign _124 = \p[124] ;
    assign _125 = \p[125] ;
    assign _126 = \p[126] ;
    assign _127 = \p[127] ;
    assign _128 = \p[128] ;
    assign _129 = \p[129] ;
    assign _130 = \p[130] ;
    assign _131 = \p[131] ;
    assign _132 = \p[132] ;
    assign _133 = \p[133] ;
    assign _134 = \p[134] ;
    assign _135 = \p[135] ;
    assign _136 = \p[136] ;
    assign _137 = \p[137] ;
    assign _138 = \p[138] ;
    assign _139 = \p[139] ;
    assign _140 = \p[140] ;
    assign _141 = \p[141] ;
    assign _142 = \p[142] ;
    assign _143 = \p[143] ;
    assign _144 = \p[144] ;
    assign _145 = \p[145] ;
    assign _146 = \p[146] ;
    assign _147 = \p[147] ;
    assign _148 = \p[148] ;
    assign _149 = \p[149] ;
    assign _150 = \p[150] ;
    assign _151 = \p[151] ;
    assign _152 = \p[152] ;
    assign _153 = \p[153] ;
    assign _154 = \p[154] ;
    assign _155 = \p[155] ;
    assign _156 = \p[156] ;
    assign _157 = \p[157] ;
    assign _158 = \p[158] ;
    assign _159 = \p[159] ;
    assign _160 = \p[160] ;
    assign _161 = \p[161] ;
    assign _162 = \p[162] ;
    assign _163 = \p[163] ;
    assign _164 = \p[164] ;
    assign _165 = \p[165] ;
    assign _166 = \p[166] ;
    assign _167 = \p[167] ;
    assign _168 = \p[168] ;
    assign _169 = \p[169] ;
    assign _170 = \p[170] ;
    assign _171 = \p[171] ;
    assign _172 = \p[172] ;
    assign _173 = \p[173] ;
    assign _174 = \p[174] ;
    assign _175 = \p[175] ;
    assign _176 = \p[176] ;
    assign _177 = \p[177] ;
    assign _178 = \p[178] ;
    assign _179 = \p[179] ;
    assign _180 = \p[180] ;
    assign _181 = \p[181] ;
    assign _182 = \p[182] ;
    assign _183 = \p[183] ;
    assign _184 = \p[184] ;
    assign _185 = \p[185] ;
    assign _186 = \p[186] ;
    assign _187 = \p[187] ;
    assign _188 = \p[188] ;
    assign _189 = \p[189] ;
    assign _190 = \p[190] ;
    assign _191 = \p[191] ;
    assign _192 = \p[192] ;
    assign _193 = \p[193] ;
    assign _194 = \p[194] ;
    assign _195 = \p[195] ;
    assign _196 = \p[196] ;
    assign _197 = \p[197] ;
    assign _198 = \p[198] ;
    assign _199 = \p[199] ;
    assign _200 = \p[200] ;
    assign _201 = \p[201] ;
    assign _202 = \p[202] ;
    assign _203 = \p[203] ;
    assign _204 = \p[204] ;
    assign _205 = \p[205] ;
    assign _206 = \p[206] ;
    assign _207 = \p[207] ;
    assign _208 = \p[208] ;
    assign _209 = \p[209] ;
    assign _210 = \p[210] ;
    assign _211 = \p[211] ;
    assign _212 = \p[212] ;
    assign _213 = \p[213] ;
    assign _214 = \p[214] ;
    assign _215 = \p[215] ;
    assign _216 = \p[216] ;
    assign _217 = \p[217] ;
    assign _218 = \p[218] ;
    assign _219 = \p[219] ;
    assign _220 = \p[220] ;
    assign _221 = \p[221] ;
    assign _222 = \p[222] ;
    assign _223 = \p[223] ;
    assign _224 = \p[224] ;
    assign _225 = \p[225] ;
    assign _226 = \p[226] ;
    assign _227 = \p[227] ;
    assign _228 = \p[228] ;
    assign _229 = \p[229] ;
    assign _230 = \p[230] ;
    assign _231 = \p[231] ;
    assign _232 = \p[232] ;
    assign _233 = \p[233] ;
    assign _234 = \p[234] ;
    assign _235 = \p[235] ;
    assign _236 = \p[236] ;
    assign _237 = \p[237] ;
    assign _238 = \p[238] ;
    assign _239 = \p[239] ;
    assign _240 = \p[240] ;
    assign _241 = \p[241] ;
    assign _242 = \p[242] ;
    assign _243 = \p[243] ;
    assign _244 = \p[244] ;
    assign _245 = \p[245] ;
    assign _246 = \p[246] ;
    assign _247 = \p[247] ;
    assign _248 = \p[248] ;
    assign _249 = \p[249] ;
    assign _250 = \p[250] ;
    assign _251 = \p[251] ;
    assign _252 = \p[252] ;
    assign _253 = \p[253] ;
    assign _254 = \p[254] ;
    assign _255 = \p[255] ;
    assign _256 = \v[0] ;
    assign _257 = \v[1] ;
    assign _258 = \v[2] ;
    assign _259 = \v[3] ;
    assign _260 = \v[4] ;
    assign _261 = \v[5] ;
    assign _262 = \v[6] ;
    assign _263 = \v[7] ;
    assign _264 = \v[8] ;
    assign _265 = \v[9] ;
    assign _266 = \v[10] ;
    assign _267 = \v[11] ;
    assign _268 = \v[12] ;
    assign _269 = \v[13] ;
    assign _270 = \v[14] ;
    assign _271 = \v[15] ;
    assign _272 = \v[16] ;
    assign _273 = \v[17] ;
    assign _274 = \v[18] ;
    assign _275 = \v[19] ;
    assign _276 = \v[20] ;
    assign _277 = \v[21] ;
    assign _278 = \v[22] ;
    assign _279 = \v[23] ;
    assign _280 = \v[24] ;
    assign _281 = \v[25] ;
    assign _282 = \v[26] ;
    assign _283 = \v[27] ;
    assign _284 = \v[28] ;
    assign _285 = \v[29] ;
    assign _286 = \v[30] ;
    assign _287 = \v[31] ;
    assign _288 = \v[32] ;
    assign _289 = \v[33] ;
    assign _290 = \v[34] ;
    assign _291 = \v[35] ;
    assign _292 = \v[36] ;
    assign _293 = \v[37] ;
    assign _294 = \v[38] ;
    assign _295 = \v[39] ;
    assign _296 = \v[40] ;
    assign _297 = \v[41] ;
    assign _298 = \v[42] ;
    assign _299 = \v[43] ;
    assign _300 = \v[44] ;
    assign _301 = \v[45] ;
    assign _302 = \v[46] ;
    assign _303 = \v[47] ;
    assign _304 = \v[48] ;
    assign _305 = \v[49] ;
    assign _306 = \v[50] ;
    assign _307 = \v[51] ;
    assign _308 = \v[52] ;
    assign _309 = \v[53] ;
    assign _310 = \v[54] ;
    assign _311 = \v[55] ;
    assign _312 = \v[56] ;
    assign _313 = \v[57] ;
    assign _314 = \v[58] ;
    assign _315 = \v[59] ;
    assign _316 = \v[60] ;
    assign _317 = \v[61] ;
    assign _318 = \v[62] ;
    assign _319 = \v[63] ;
    assign _320 = \v[64] ;
    assign _321 = \v[65] ;
    assign _322 = \v[66] ;
    assign _323 = \v[67] ;
    assign _324 = \v[68] ;
    assign _325 = \v[69] ;
    assign _326 = \v[70] ;
    assign _327 = \v[71] ;
    assign _328 = \v[72] ;
    assign _329 = \v[73] ;
    assign _330 = \v[74] ;
    assign _331 = \v[75] ;
    assign _332 = \v[76] ;
    assign _333 = \v[77] ;
    assign _334 = \v[78] ;
    assign _335 = \v[79] ;
    assign _336 = \v[80] ;
    assign _337 = \v[81] ;
    assign _338 = \v[82] ;
    assign _339 = \v[83] ;
    assign _340 = \v[84] ;
    assign _341 = \v[85] ;
    assign _342 = \v[86] ;
    assign _343 = \v[87] ;
    assign _344 = \v[88] ;
    assign _345 = \v[89] ;
    assign _346 = \v[90] ;
    assign _347 = \v[91] ;
    assign _348 = \v[92] ;
    assign _349 = \v[93] ;
    assign _350 = \v[94] ;
    assign _351 = \v[95] ;
    assign _352 = \v[96] ;
    assign _353 = \v[97] ;
    assign _354 = \v[98] ;
    assign _355 = \v[99] ;
    assign _356 = \v[100] ;
    assign _357 = \v[101] ;
    assign _358 = \v[102] ;
    assign _359 = \v[103] ;
    assign _360 = \v[104] ;
    assign _361 = \v[105] ;
    assign _362 = \v[106] ;
    assign _363 = \v[107] ;
    assign _364 = \v[108] ;
    assign _365 = \v[109] ;
    assign _366 = \v[110] ;
    assign _367 = \v[111] ;
    assign _368 = \v[112] ;
    assign _369 = \v[113] ;
    assign _370 = \v[114] ;
    assign _371 = \v[115] ;
    assign _372 = \v[116] ;
    assign _373 = \v[117] ;
    assign _374 = \v[118] ;
    assign _375 = \v[119] ;
    assign _376 = \v[120] ;
    assign _377 = \v[121] ;
    assign _378 = \v[122] ;
    assign _379 = \v[123] ;
    assign _380 = \v[124] ;
    assign _381 = \v[125] ;
    assign _382 = \v[126] ;
    assign _383 = \v[127] ;
    assign _384 = \v[128] ;
    assign _385 = \v[129] ;
    assign _386 = \v[130] ;
    assign _387 = \v[131] ;
    assign _388 = \v[132] ;
    assign _389 = \v[133] ;
    assign _390 = \v[134] ;
    assign _391 = \v[135] ;
    assign _392 = \v[136] ;
    assign _393 = \v[137] ;
    assign _394 = \v[138] ;
    assign _395 = \v[139] ;
    assign _396 = \v[140] ;
    assign _397 = \v[141] ;
    assign _398 = \v[142] ;
    assign _399 = \v[143] ;
    assign _400 = \v[144] ;
    assign _401 = \v[145] ;
    assign _402 = \v[146] ;
    assign _403 = \v[147] ;
    assign _404 = \v[148] ;
    assign _405 = \v[149] ;
    assign _406 = \v[150] ;
    assign _407 = \v[151] ;
    assign _408 = \v[152] ;
    assign _409 = \v[153] ;
    assign _410 = \v[154] ;
    assign _411 = \v[155] ;
    assign _412 = \v[156] ;
    assign _413 = \v[157] ;
    assign _414 = \v[158] ;
    assign _415 = \v[159] ;
    assign _416 = \v[160] ;
    assign _417 = \v[161] ;
    assign _418 = \v[162] ;
    assign _419 = \v[163] ;
    assign _420 = \v[164] ;
    assign _421 = \v[165] ;
    assign _422 = \v[166] ;
    assign _423 = \v[167] ;
    assign _424 = \v[168] ;
    assign _425 = \v[169] ;
    assign _426 = \v[170] ;
    assign _427 = \v[171] ;
    assign _428 = \v[172] ;
    assign _429 = \v[173] ;
    assign _430 = \v[174] ;
    assign _431 = \v[175] ;
    assign _432 = \v[176] ;
    assign _433 = \v[177] ;
    assign _434 = \v[178] ;
    assign _435 = \v[179] ;
    assign _436 = \v[180] ;
    assign _437 = \v[181] ;
    assign _438 = \v[182] ;
    assign _439 = \v[183] ;
    assign _440 = \v[184] ;
    assign _441 = \v[185] ;
    assign _442 = \v[186] ;
    assign _443 = \v[187] ;
    assign _444 = \v[188] ;
    assign _445 = \v[189] ;
    assign _446 = \v[190] ;
    assign _447 = \v[191] ;
    assign _448 = \v[192] ;
    assign _449 = \v[193] ;
    assign _450 = \v[194] ;
    assign _451 = \v[195] ;
    assign _452 = \v[196] ;
    assign _453 = \v[197] ;
    assign _454 = \v[198] ;
    assign _455 = \v[199] ;
    assign _456 = \v[200] ;
    assign _457 = \v[201] ;
    assign _458 = \v[202] ;
    assign _459 = \v[203] ;
    assign _460 = \v[204] ;
    assign _461 = \v[205] ;
    assign _462 = \v[206] ;
    assign _463 = \v[207] ;
    assign _464 = \v[208] ;
    assign _465 = \v[209] ;
    assign _466 = \v[210] ;
    assign _467 = \v[211] ;
    assign _468 = \v[212] ;
    assign _469 = \v[213] ;
    assign _470 = \v[214] ;
    assign _471 = \v[215] ;
    assign _472 = \v[216] ;
    assign _473 = \v[217] ;
    assign _474 = \v[218] ;
    assign _475 = \v[219] ;
    assign _476 = \v[220] ;
    assign _477 = \v[221] ;
    assign _478 = \v[222] ;
    assign _479 = \v[223] ;
    assign _480 = \v[224] ;
    assign _481 = \v[225] ;
    assign _482 = \v[226] ;
    assign _483 = \v[227] ;
    assign _484 = \v[228] ;
    assign _485 = \v[229] ;
    assign _486 = \v[230] ;
    assign _487 = \v[231] ;
    assign _488 = \v[232] ;
    assign _489 = \v[233] ;
    assign _490 = \v[234] ;
    assign _491 = \v[235] ;
    assign _492 = \v[236] ;
    assign _493 = \v[237] ;
    assign _494 = \v[238] ;
    assign _495 = \v[239] ;
    assign _496 = \v[240] ;
    assign _497 = \v[241] ;
    assign _498 = \v[242] ;
    assign _499 = \v[243] ;
    assign _500 = \v[244] ;
    assign _501 = \v[245] ;
    assign _502 = \v[246] ;
    assign _503 = \v[247] ;
    assign _504 = \v[248] ;
    assign _505 = \v[249] ;
    assign _506 = \v[250] ;
    assign _507 = \v[251] ;
    assign _508 = \v[252] ;
    assign _509 = \v[253] ;
    assign _510 = \v[254] ;
    assign _511 = \v[255] ;
    assign _512 = _0 | _1;
    assign _513 = _0 & _256;
    assign _514 = !_0;
    assign _515 = _514 & _257;
    assign _516 = _513 | _515;
    assign _517 = _2 | _3;
    assign _518 = _2 & _258;
    assign _519 = !_2;
    assign _520 = _519 & _259;
    assign _521 = _518 | _520;
    assign _522 = _512 | _517;
    assign _523 = _512 & _516;
    assign _524 = !_512;
    assign _525 = _524 & _521;
    assign _526 = _523 | _525;
    assign _527 = _4 | _5;
    assign _528 = _4 & _260;
    assign _529 = !_4;
    assign _530 = _529 & _261;
    assign _531 = _528 | _530;
    assign _532 = _6 | _7;
    assign _533 = _6 & _262;
    assign _534 = !_6;
    assign _535 = _534 & _263;
    assign _536 = _533 | _535;
    assign _537 = _527 | _532;
    assign _538 = _527 & _531;
    assign _539 = !_527;
    assign _540 = _539 & _536;
    assign _541 = _538 | _540;
    assign _542 = _522 | _537;
    assign _543 = _522 & _526;
    assign _544 = !_522;
    assign _545 = _544 & _541;
    assign _546 = _543 | _545;
    assign _547 = _8 | _9;
    assign _548 = _8 & _264;
    assign _549 = !_8;
    assign _550 = _549 & _265;
    assign _551 = _548 | _550;
    assign _552 = _10 | _11;
    assign _553 = _10 & _266;
    assign _554 = !_10;
    assign _555 = _554 & _267;
    assign _556 = _553 | _555;
    assign _557 = _547 | _552;
    assign _558 = _547 & _551;
    assign _559 = !_547;
    assign _560 = _559 & _556;
    assign _561 = _558 | _560;
    assign _562 = _12 | _13;
    assign _563 = _12 & _268;
    assign _564 = !_12;
    assign _565 = _564 & _269;
    assign _566 = _563 | _565;
    assign _567 = _14 | _15;
    assign _568 = _14 & _270;
    assign _569 = !_14;
    assign _570 = _569 & _271;
    assign _571 = _568 | _570;
    assign _572 = _562 | _567;
    assign _573 = _562 & _566;
    assign _574 = !_562;
    assign _575 = _574 & _571;
    assign _576 = _573 | _575;
    assign _577 = _557 | _572;
    assign _578 = _557 & _561;
    assign _579 = !_557;
    assign _580 = _579 & _576;
    assign _581 = _578 | _580;
    assign _582 = _542 | _577;
    assign _583 = _542 & _546;
    assign _584 = !_542;
    assign _585 = _584 & _581;
    assign _586 = _583 | _585;
    assign _587 = _16 | _17;
    assign _588 = _16 & _272;
    assign _589 = !_16;
    assign _590 = _589 & _273;
    assign _591 = _588 | _590;
    assign _592 = _18 | _19;
    assign _593 = _18 & _274;
    assign _594 = !_18;
    assign _595 = _594 & _275;
    assign _596 = _593 | _595;
    assign _597 = _587 | _592;
    assign _598 = _587 & _591;
    assign _599 = !_587;
    assign _600 = _599 & _596;
    assign _601 = _598 | _600;
    assign _602 = _20 | _21;
    assign _603 = _20 & _276;
    assign _604 = !_20;
    assign _605 = _604 & _277;
    assign _606 = _603 | _605;
    assign _607 = _22 | _23;
    assign _608 = _22 & _278;
    assign _609 = !_22;
    assign _610 = _609 & _279;
    assign _611 = _608 | _610;
    assign _612 = _602 | _607;
    assign _613 = _602 & _606;
    assign _614 = !_602;
    assign _615 = _614 & _611;
    assign _616 = _613 | _615;
    assign _617 = _597 | _612;
    assign _618 = _597 & _601;
    assign _619 = !_597;
    assign _620 = _619 & _616;
    assign _621 = _618 | _620;
    assign _622 = _24 | _25;
    assign _623 = _24 & _280;
    assign _624 = !_24;
    assign _625 = _624 & _281;
    assign _626 = _623 | _625;
    assign _627 = _26 | _27;
    assign _628 = _26 & _282;
    assign _629 = !_26;
    assign _630 = _629 & _283;
    assign _631 = _628 | _630;
    assign _632 = _622 | _627;
    assign _633 = _622 & _626;
    assign _634 = !_622;
    assign _635 = _634 & _631;
    assign _636 = _633 | _635;
    assign _637 = _28 | _29;
    assign _638 = _28 & _284;
    assign _639 = !_28;
    assign _640 = _639 & _285;
    assign _641 = _638 | _640;
    assign _642 = _30 | _31;
    assign _643 = _30 & _286;
    assign _644 = !_30;
    assign _645 = _644 & _287;
    assign _646 = _643 | _645;
    assign _647 = _637 | _642;
    assign _648 = _637 & _641;
    assign _649 = !_637;
    assign _650 = _649 & _646;
    assign _651 = _648 | _650;
    assign _652 = _632 | _647;
    assign _653 = _632 & _636;
    assign _654 = !_632;
    assign _655 = _654 & _651;
    assign _656 = _653 | _655;
    assign _657 = _617 | _652;
    assign _658 = _617 & _621;
    assign _659 = !_617;
    assign _660 = _659 & _656;
    assign _661 = _658 | _660;
    assign _662 = _582 | _657;
    assign _663 = _582 & _586;
    assign _664 = !_582;
    assign _665 = _664 & _661;
    assign _666 = _663 | _665;
    assign _667 = _32 | _33;
    assign _668 = _32 & _288;
    assign _669 = !_32;
    assign _670 = _669 & _289;
    assign _671 = _668 | _670;
    assign _672 = _34 | _35;
    assign _673 = _34 & _290;
    assign _674 = !_34;
    assign _675 = _674 & _291;
    assign _676 = _673 | _675;
    assign _677 = _667 | _672;
    assign _678 = _667 & _671;
    assign _679 = !_667;
    assign _680 = _679 & _676;
    assign _681 = _678 | _680;
    assign _682 = _36 | _37;
    assign _683 = _36 & _292;
    assign _684 = !_36;
    assign _685 = _684 & _293;
    assign _686 = _683 | _685;
    assign _687 = _38 | _39;
    assign _688 = _38 & _294;
    assign _689 = !_38;
    assign _690 = _689 & _295;
    assign _691 = _688 | _690;
    assign _692 = _682 | _687;
    assign _693 = _682 & _686;
    assign _694 = !_682;
    assign _695 = _694 & _691;
    assign _696 = _693 | _695;
    assign _697 = _677 | _692;
    assign _698 = _677 & _681;
    assign _699 = !_677;
    assign _700 = _699 & _696;
    assign _701 = _698 | _700;
    assign _702 = _40 | _41;
    assign _703 = _40 & _296;
    assign _704 = !_40;
    assign _705 = _704 & _297;
    assign _706 = _703 | _705;
    assign _707 = _42 | _43;
    assign _708 = _42 & _298;
    assign _709 = !_42;
    assign _710 = _709 & _299;
    assign _711 = _708 | _710;
    assign _712 = _702 | _707;
    assign _713 = _702 & _706;
    assign _714 = !_702;
    assign _715 = _714 & _711;
    assign _716 = _713 | _715;
    assign _717 = _44 | _45;
    assign _718 = _44 & _300;
    assign _719 = !_44;
    assign _720 = _719 & _301;
    assign _721 = _718 | _720;
    assign _722 = _46 | _47;
    assign _723 = _46 & _302;
    assign _724 = !_46;
    assign _725 = _724 & _303;
    assign _726 = _723 | _725;
    assign _727 = _717 | _722;
    assign _728 = _717 & _721;
    assign _729 = !_717;
    assign _730 = _729 & _726;
    assign _731 = _728 | _730;
    assign _732 = _712 | _727;
    assign _733 = _712 & _716;
    assign _734 = !_712;
    assign _735 = _734 & _731;
    assign _736 = _733 | _735;
    assign _737 = _697 | _732;
    assign _738 = _697 & _701;
    assign _739 = !_697;
    assign _740 = _739 & _736;
    assign _741 = _738 | _740;
    assign _742 = _48 | _49;
    assign _743 = _48 & _304;
    assign _744 = !_48;
    assign _745 = _744 & _305;
    assign _746 = _743 | _745;
    assign _747 = _50 | _51;
    assign _748 = _50 & _306;
    assign _749 = !_50;
    assign _750 = _749 & _307;
    assign _751 = _748 | _750;
    assign _752 = _742 | _747;
    assign _753 = _742 & _746;
    assign _754 = !_742;
    assign _755 = _754 & _751;
    assign _756 = _753 | _755;
    assign _757 = _52 | _53;
    assign _758 = _52 & _308;
    assign _759 = !_52;
    assign _760 = _759 & _309;
    assign _761 = _758 | _760;
    assign _762 = _54 | _55;
    assign _763 = _54 & _310;
    assign _764 = !_54;
    assign _765 = _764 & _311;
    assign _766 = _763 | _765;
    assign _767 = _757 | _762;
    assign _768 = _757 & _761;
    assign _769 = !_757;
    assign _770 = _769 & _766;
    assign _771 = _768 | _770;
    assign _772 = _752 | _767;
    assign _773 = _752 & _756;
    assign _774 = !_752;
    assign _775 = _774 & _771;
    assign _776 = _773 | _775;
    assign _777 = _56 | _57;
    assign _778 = _56 & _312;
    assign _779 = !_56;
    assign _780 = _779 & _313;
    assign _781 = _778 | _780;
    assign _782 = _58 | _59;
    assign _783 = _58 & _314;
    assign _784 = !_58;
    assign _785 = _784 & _315;
    assign _786 = _783 | _785;
    assign _787 = _777 | _782;
    assign _788 = _777 & _781;
    assign _789 = !_777;
    assign _790 = _789 & _786;
    assign _791 = _788 | _790;
    assign _792 = _60 | _61;
    assign _793 = _60 & _316;
    assign _794 = !_60;
    assign _795 = _794 & _317;
    assign _796 = _793 | _795;
    assign _797 = _62 | _63;
    assign _798 = _62 & _318;
    assign _799 = !_62;
    assign _800 = _799 & _319;
    assign _801 = _798 | _800;
    assign _802 = _792 | _797;
    assign _803 = _792 & _796;
    assign _804 = !_792;
    assign _805 = _804 & _801;
    assign _806 = _803 | _805;
    assign _807 = _787 | _802;
    assign _808 = _787 & _791;
    assign _809 = !_787;
    assign _810 = _809 & _806;
    assign _811 = _808 | _810;
    assign _812 = _772 | _807;
    assign _813 = _772 & _776;
    assign _814 = !_772;
    assign _815 = _814 & _811;
    assign _816 = _813 | _815;
    assign _817 = _737 | _812;
    assign _818 = _737 & _741;
    assign _819 = !_737;
    assign _820 = _819 & _816;
    assign _821 = _818 | _820;
    assign _822 = _662 | _817;
    assign _823 = _662 & _666;
    assign _824 = !_662;
    assign _825 = _824 & _821;
    assign _826 = _823 | _825;
    assign _827 = _64 | _65;
    assign _828 = _64 & _320;
    assign _829 = !_64;
    assign _830 = _829 & _321;
    assign _831 = _828 | _830;
    assign _832 = _66 | _67;
    assign _833 = _66 & _322;
    assign _834 = !_66;
    assign _835 = _834 & _323;
    assign _836 = _833 | _835;
    assign _837 = _827 | _832;
    assign _838 = _827 & _831;
    assign _839 = !_827;
    assign _840 = _839 & _836;
    assign _841 = _838 | _840;
    assign _842 = _68 | _69;
    assign _843 = _68 & _324;
    assign _844 = !_68;
    assign _845 = _844 & _325;
    assign _846 = _843 | _845;
    assign _847 = _70 | _71;
    assign _848 = _70 & _326;
    assign _849 = !_70;
    assign _850 = _849 & _327;
    assign _851 = _848 | _850;
    assign _852 = _842 | _847;
    assign _853 = _842 & _846;
    assign _854 = !_842;
    assign _855 = _854 & _851;
    assign _856 = _853 | _855;
    assign _857 = _837 | _852;
    assign _858 = _837 & _841;
    assign _859 = !_837;
    assign _860 = _859 & _856;
    assign _861 = _858 | _860;
    assign _862 = _72 | _73;
    assign _863 = _72 & _328;
    assign _864 = !_72;
    assign _865 = _864 & _329;
    assign _866 = _863 | _865;
    assign _867 = _74 | _75;
    assign _868 = _74 & _330;
    assign _869 = !_74;
    assign _870 = _869 & _331;
    assign _871 = _868 | _870;
    assign _872 = _862 | _867;
    assign _873 = _862 & _866;
    assign _874 = !_862;
    assign _875 = _874 & _871;
    assign _876 = _873 | _875;
    assign _877 = _76 | _77;
    assign _878 = _76 & _332;
    assign _879 = !_76;
    assign _880 = _879 & _333;
    assign _881 = _878 | _880;
    assign _882 = _78 | _79;
    assign _883 = _78 & _334;
    assign _884 = !_78;
    assign _885 = _884 & _335;
    assign _886 = _883 | _885;
    assign _887 = _877 | _882;
    assign _888 = _877 & _881;
    assign _889 = !_877;
    assign _890 = _889 & _886;
    assign _891 = _888 | _890;
    assign _892 = _872 | _887;
    assign _893 = _872 & _876;
    assign _894 = !_872;
    assign _895 = _894 & _891;
    assign _896 = _893 | _895;
    assign _897 = _857 | _892;
    assign _898 = _857 & _861;
    assign _899 = !_857;
    assign _900 = _899 & _896;
    assign _901 = _898 | _900;
    assign _902 = _80 | _81;
    assign _903 = _80 & _336;
    assign _904 = !_80;
    assign _905 = _904 & _337;
    assign _906 = _903 | _905;
    assign _907 = _82 | _83;
    assign _908 = _82 & _338;
    assign _909 = !_82;
    assign _910 = _909 & _339;
    assign _911 = _908 | _910;
    assign _912 = _902 | _907;
    assign _913 = _902 & _906;
    assign _914 = !_902;
    assign _915 = _914 & _911;
    assign _916 = _913 | _915;
    assign _917 = _84 | _85;
    assign _918 = _84 & _340;
    assign _919 = !_84;
    assign _920 = _919 & _341;
    assign _921 = _918 | _920;
    assign _922 = _86 | _87;
    assign _923 = _86 & _342;
    assign _924 = !_86;
    assign _925 = _924 & _343;
    assign _926 = _923 | _925;
    assign _927 = _917 | _922;
    assign _928 = _917 & _921;
    assign _929 = !_917;
    assign _930 = _929 & _926;
    assign _931 = _928 | _930;
    assign _932 = _912 | _927;
    assign _933 = _912 & _916;
    assign _934 = !_912;
    assign _935 = _934 & _931;
    assign _936 = _933 | _935;
    assign _937 = _88 | _89;
    assign _938 = _88 & _344;
    assign _939 = !_88;
    assign _940 = _939 & _345;
    assign _941 = _938 | _940;
    assign _942 = _90 | _91;
    assign _943 = _90 & _346;
    assign _944 = !_90;
    assign _945 = _944 & _347;
    assign _946 = _943 | _945;
    assign _947 = _937 | _942;
    assign _948 = _937 & _941;
    assign _949 = !_937;
    assign _950 = _949 & _946;
    assign _951 = _948 | _950;
    assign _952 = _92 | _93;
    assign _953 = _92 & _348;
    assign _954 = !_92;
    assign _955 = _954 & _349;
    assign _956 = _953 | _955;
    assign _957 = _94 | _95;
    assign _958 = _94 & _350;
    assign _959 = !_94;
    assign _960 = _959 & _351;
    assign _961 = _958 | _960;
    assign _962 = _952 | _957;
    assign _963 = _952 & _956;
    assign _964 = !_952;
    assign _965 = _964 & _961;
    assign _966 = _963 | _965;
    assign _967 = _947 | _962;
    assign _968 = _947 & _951;
    assign _969 = !_947;
    assign _970 = _969 & _966;
    assign _971 = _968 | _970;
    assign _972 = _932 | _967;
    assign _973 = _932 & _936;
    assign _974 = !_932;
    assign _975 = _974 & _971;
    assign _976 = _973 | _975;
    assign _977 = _897 | _972;
    assign _978 = _897 & _901;
    assign _979 = !_897;
    assign _980 = _979 & _976;
    assign _981 = _978 | _980;
    assign _982 = _96 | _97;
    assign _983 = _96 & _352;
    assign _984 = !_96;
    assign _985 = _984 & _353;
    assign _986 = _983 | _985;
    assign _987 = _98 | _99;
    assign _988 = _98 & _354;
    assign _989 = !_98;
    assign _990 = _989 & _355;
    assign _991 = _988 | _990;
    assign _992 = _982 | _987;
    assign _993 = _982 & _986;
    assign _994 = !_982;
    assign _995 = _994 & _991;
    assign _996 = _993 | _995;
    assign _997 = _100 | _101;
    assign _998 = _100 & _356;
    assign _999 = !_100;
    assign _1000 = _999 & _357;
    assign _1001 = _998 | _1000;
    assign _1002 = _102 | _103;
    assign _1003 = _102 & _358;
    assign _1004 = !_102;
    assign _1005 = _1004 & _359;
    assign _1006 = _1003 | _1005;
    assign _1007 = _997 | _1002;
    assign _1008 = _997 & _1001;
    assign _1009 = !_997;
    assign _1010 = _1009 & _1006;
    assign _1011 = _1008 | _1010;
    assign _1012 = _992 | _1007;
    assign _1013 = _992 & _996;
    assign _1014 = !_992;
    assign _1015 = _1014 & _1011;
    assign _1016 = _1013 | _1015;
    assign _1017 = _104 | _105;
    assign _1018 = _104 & _360;
    assign _1019 = !_104;
    assign _1020 = _1019 & _361;
    assign _1021 = _1018 | _1020;
    assign _1022 = _106 | _107;
    assign _1023 = _106 & _362;
    assign _1024 = !_106;
    assign _1025 = _1024 & _363;
    assign _1026 = _1023 | _1025;
    assign _1027 = _1017 | _1022;
    assign _1028 = _1017 & _1021;
    assign _1029 = !_1017;
    assign _1030 = _1029 & _1026;
    assign _1031 = _1028 | _1030;
    assign _1032 = _108 | _109;
    assign _1033 = _108 & _364;
    assign _1034 = !_108;
    assign _1035 = _1034 & _365;
    assign _1036 = _1033 | _1035;
    assign _1037 = _110 | _111;
    assign _1038 = _110 & _366;
    assign _1039 = !_110;
    assign _1040 = _1039 & _367;
    assign _1041 = _1038 | _1040;
    assign _1042 = _1032 | _1037;
    assign _1043 = _1032 & _1036;
    assign _1044 = !_1032;
    assign _1045 = _1044 & _1041;
    assign _1046 = _1043 | _1045;
    assign _1047 = _1027 | _1042;
    assign _1048 = _1027 & _1031;
    assign _1049 = !_1027;
    assign _1050 = _1049 & _1046;
    assign _1051 = _1048 | _1050;
    assign _1052 = _1012 | _1047;
    assign _1053 = _1012 & _1016;
    assign _1054 = !_1012;
    assign _1055 = _1054 & _1051;
    assign _1056 = _1053 | _1055;
    assign _1057 = _112 | _113;
    assign _1058 = _112 & _368;
    assign _1059 = !_112;
    assign _1060 = _1059 & _369;
    assign _1061 = _1058 | _1060;
    assign _1062 = _114 | _115;
    assign _1063 = _114 & _370;
    assign _1064 = !_114;
    assign _1065 = _1064 & _371;
    assign _1066 = _1063 | _1065;
    assign _1067 = _1057 | _1062;
    assign _1068 = _1057 & _1061;
    assign _1069 = !_1057;
    assign _1070 = _1069 & _1066;
    assign _1071 = _1068 | _1070;
    assign _1072 = _116 | _117;
    assign _1073 = _116 & _372;
    assign _1074 = !_116;
    assign _1075 = _1074 & _373;
    assign _1076 = _1073 | _1075;
    assign _1077 = _118 | _119;
    assign _1078 = _118 & _374;
    assign _1079 = !_118;
    assign _1080 = _1079 & _375;
    assign _1081 = _1078 | _1080;
    assign _1082 = _1072 | _1077;
    assign _1083 = _1072 & _1076;
    assign _1084 = !_1072;
    assign _1085 = _1084 & _1081;
    assign _1086 = _1083 | _1085;
    assign _1087 = _1067 | _1082;
    assign _1088 = _1067 & _1071;
    assign _1089 = !_1067;
    assign _1090 = _1089 & _1086;
    assign _1091 = _1088 | _1090;
    assign _1092 = _120 | _121;
    assign _1093 = _120 & _376;
    assign _1094 = !_120;
    assign _1095 = _1094 & _377;
    assign _1096 = _1093 | _1095;
    assign _1097 = _122 | _123;
    assign _1098 = _122 & _378;
    assign _1099 = !_122;
    assign _1100 = _1099 & _379;
    assign _1101 = _1098 | _1100;
    assign _1102 = _1092 | _1097;
    assign _1103 = _1092 & _1096;
    assign _1104 = !_1092;
    assign _1105 = _1104 & _1101;
    assign _1106 = _1103 | _1105;
    assign _1107 = _124 | _125;
    assign _1108 = _124 & _380;
    assign _1109 = !_124;
    assign _1110 = _1109 & _381;
    assign _1111 = _1108 | _1110;
    assign _1112 = _126 | _127;
    assign _1113 = _126 & _382;
    assign _1114 = !_126;
    assign _1115 = _1114 & _383;
    assign _1116 = _1113 | _1115;
    assign _1117 = _1107 | _1112;
    assign _1118 = _1107 & _1111;
    assign _1119 = !_1107;
    assign _1120 = _1119 & _1116;
    assign _1121 = _1118 | _1120;
    assign _1122 = _1102 | _1117;
    assign _1123 = _1102 & _1106;
    assign _1124 = !_1102;
    assign _1125 = _1124 & _1121;
    assign _1126 = _1123 | _1125;
    assign _1127 = _1087 | _1122;
    assign _1128 = _1087 & _1091;
    assign _1129 = !_1087;
    assign _1130 = _1129 & _1126;
    assign _1131 = _1128 | _1130;
    assign _1132 = _1052 | _1127;
    assign _1133 = _1052 & _1056;
    assign _1134 = !_1052;
    assign _1135 = _1134 & _1131;
    assign _1136 = _1133 | _1135;
    assign _1137 = _977 | _1132;
    assign _1138 = _977 & _981;
    assign _1139 = !_977;
    assign _1140 = _1139 & _1136;
    assign _1141 = _1138 | _1140;
    assign _1142 = _822 | _1137;
    assign _1143 = _822 & _826;
    assign _1144 = !_822;
    assign _1145 = _1144 & _1141;
    assign _1146 = _1143 | _1145;
    assign _1147 = _128 | _129;
    assign _1148 = _128 & _384;
    assign _1149 = !_128;
    assign _1150 = _1149 & _385;
    assign _1151 = _1148 | _1150;
    assign _1152 = _130 | _131;
    assign _1153 = _130 & _386;
    assign _1154 = !_130;
    assign _1155 = _1154 & _387;
    assign _1156 = _1153 | _1155;
    assign _1157 = _1147 | _1152;
    assign _1158 = _1147 & _1151;
    assign _1159 = !_1147;
    assign _1160 = _1159 & _1156;
    assign _1161 = _1158 | _1160;
    assign _1162 = _132 | _133;
    assign _1163 = _132 & _388;
    assign _1164 = !_132;
    assign _1165 = _1164 & _389;
    assign _1166 = _1163 | _1165;
    assign _1167 = _134 | _135;
    assign _1168 = _134 & _390;
    assign _1169 = !_134;
    assign _1170 = _1169 & _391;
    assign _1171 = _1168 | _1170;
    assign _1172 = _1162 | _1167;
    assign _1173 = _1162 & _1166;
    assign _1174 = !_1162;
    assign _1175 = _1174 & _1171;
    assign _1176 = _1173 | _1175;
    assign _1177 = _1157 | _1172;
    assign _1178 = _1157 & _1161;
    assign _1179 = !_1157;
    assign _1180 = _1179 & _1176;
    assign _1181 = _1178 | _1180;
    assign _1182 = _136 | _137;
    assign _1183 = _136 & _392;
    assign _1184 = !_136;
    assign _1185 = _1184 & _393;
    assign _1186 = _1183 | _1185;
    assign _1187 = _138 | _139;
    assign _1188 = _138 & _394;
    assign _1189 = !_138;
    assign _1190 = _1189 & _395;
    assign _1191 = _1188 | _1190;
    assign _1192 = _1182 | _1187;
    assign _1193 = _1182 & _1186;
    assign _1194 = !_1182;
    assign _1195 = _1194 & _1191;
    assign _1196 = _1193 | _1195;
    assign _1197 = _140 | _141;
    assign _1198 = _140 & _396;
    assign _1199 = !_140;
    assign _1200 = _1199 & _397;
    assign _1201 = _1198 | _1200;
    assign _1202 = _142 | _143;
    assign _1203 = _142 & _398;
    assign _1204 = !_142;
    assign _1205 = _1204 & _399;
    assign _1206 = _1203 | _1205;
    assign _1207 = _1197 | _1202;
    assign _1208 = _1197 & _1201;
    assign _1209 = !_1197;
    assign _1210 = _1209 & _1206;
    assign _1211 = _1208 | _1210;
    assign _1212 = _1192 | _1207;
    assign _1213 = _1192 & _1196;
    assign _1214 = !_1192;
    assign _1215 = _1214 & _1211;
    assign _1216 = _1213 | _1215;
    assign _1217 = _1177 | _1212;
    assign _1218 = _1177 & _1181;
    assign _1219 = !_1177;
    assign _1220 = _1219 & _1216;
    assign _1221 = _1218 | _1220;
    assign _1222 = _144 | _145;
    assign _1223 = _144 & _400;
    assign _1224 = !_144;
    assign _1225 = _1224 & _401;
    assign _1226 = _1223 | _1225;
    assign _1227 = _146 | _147;
    assign _1228 = _146 & _402;
    assign _1229 = !_146;
    assign _1230 = _1229 & _403;
    assign _1231 = _1228 | _1230;
    assign _1232 = _1222 | _1227;
    assign _1233 = _1222 & _1226;
    assign _1234 = !_1222;
    assign _1235 = _1234 & _1231;
    assign _1236 = _1233 | _1235;
    assign _1237 = _148 | _149;
    assign _1238 = _148 & _404;
    assign _1239 = !_148;
    assign _1240 = _1239 & _405;
    assign _1241 = _1238 | _1240;
    assign _1242 = _150 | _151;
    assign _1243 = _150 & _406;
    assign _1244 = !_150;
    assign _1245 = _1244 & _407;
    assign _1246 = _1243 | _1245;
    assign _1247 = _1237 | _1242;
    assign _1248 = _1237 & _1241;
    assign _1249 = !_1237;
    assign _1250 = _1249 & _1246;
    assign _1251 = _1248 | _1250;
    assign _1252 = _1232 | _1247;
    assign _1253 = _1232 & _1236;
    assign _1254 = !_1232;
    assign _1255 = _1254 & _1251;
    assign _1256 = _1253 | _1255;
    assign _1257 = _152 | _153;
    assign _1258 = _152 & _408;
    assign _1259 = !_152;
    assign _1260 = _1259 & _409;
    assign _1261 = _1258 | _1260;
    assign _1262 = _154 | _155;
    assign _1263 = _154 & _410;
    assign _1264 = !_154;
    assign _1265 = _1264 & _411;
    assign _1266 = _1263 | _1265;
    assign _1267 = _1257 | _1262;
    assign _1268 = _1257 & _1261;
    assign _1269 = !_1257;
    assign _1270 = _1269 & _1266;
    assign _1271 = _1268 | _1270;
    assign _1272 = _156 | _157;
    assign _1273 = _156 & _412;
    assign _1274 = !_156;
    assign _1275 = _1274 & _413;
    assign _1276 = _1273 | _1275;
    assign _1277 = _158 | _159;
    assign _1278 = _158 & _414;
    assign _1279 = !_158;
    assign _1280 = _1279 & _415;
    assign _1281 = _1278 | _1280;
    assign _1282 = _1272 | _1277;
    assign _1283 = _1272 & _1276;
    assign _1284 = !_1272;
    assign _1285 = _1284 & _1281;
    assign _1286 = _1283 | _1285;
    assign _1287 = _1267 | _1282;
    assign _1288 = _1267 & _1271;
    assign _1289 = !_1267;
    assign _1290 = _1289 & _1286;
    assign _1291 = _1288 | _1290;
    assign _1292 = _1252 | _1287;
    assign _1293 = _1252 & _1256;
    assign _1294 = !_1252;
    assign _1295 = _1294 & _1291;
    assign _1296 = _1293 | _1295;
    assign _1297 = _1217 | _1292;
    assign _1298 = _1217 & _1221;
    assign _1299 = !_1217;
    assign _1300 = _1299 & _1296;
    assign _1301 = _1298 | _1300;
    assign _1302 = _160 | _161;
    assign _1303 = _160 & _416;
    assign _1304 = !_160;
    assign _1305 = _1304 & _417;
    assign _1306 = _1303 | _1305;
    assign _1307 = _162 | _163;
    assign _1308 = _162 & _418;
    assign _1309 = !_162;
    assign _1310 = _1309 & _419;
    assign _1311 = _1308 | _1310;
    assign _1312 = _1302 | _1307;
    assign _1313 = _1302 & _1306;
    assign _1314 = !_1302;
    assign _1315 = _1314 & _1311;
    assign _1316 = _1313 | _1315;
    assign _1317 = _164 | _165;
    assign _1318 = _164 & _420;
    assign _1319 = !_164;
    assign _1320 = _1319 & _421;
    assign _1321 = _1318 | _1320;
    assign _1322 = _166 | _167;
    assign _1323 = _166 & _422;
    assign _1324 = !_166;
    assign _1325 = _1324 & _423;
    assign _1326 = _1323 | _1325;
    assign _1327 = _1317 | _1322;
    assign _1328 = _1317 & _1321;
    assign _1329 = !_1317;
    assign _1330 = _1329 & _1326;
    assign _1331 = _1328 | _1330;
    assign _1332 = _1312 | _1327;
    assign _1333 = _1312 & _1316;
    assign _1334 = !_1312;
    assign _1335 = _1334 & _1331;
    assign _1336 = _1333 | _1335;
    assign _1337 = _168 | _169;
    assign _1338 = _168 & _424;
    assign _1339 = !_168;
    assign _1340 = _1339 & _425;
    assign _1341 = _1338 | _1340;
    assign _1342 = _170 | _171;
    assign _1343 = _170 & _426;
    assign _1344 = !_170;
    assign _1345 = _1344 & _427;
    assign _1346 = _1343 | _1345;
    assign _1347 = _1337 | _1342;
    assign _1348 = _1337 & _1341;
    assign _1349 = !_1337;
    assign _1350 = _1349 & _1346;
    assign _1351 = _1348 | _1350;
    assign _1352 = _172 | _173;
    assign _1353 = _172 & _428;
    assign _1354 = !_172;
    assign _1355 = _1354 & _429;
    assign _1356 = _1353 | _1355;
    assign _1357 = _174 | _175;
    assign _1358 = _174 & _430;
    assign _1359 = !_174;
    assign _1360 = _1359 & _431;
    assign _1361 = _1358 | _1360;
    assign _1362 = _1352 | _1357;
    assign _1363 = _1352 & _1356;
    assign _1364 = !_1352;
    assign _1365 = _1364 & _1361;
    assign _1366 = _1363 | _1365;
    assign _1367 = _1347 | _1362;
    assign _1368 = _1347 & _1351;
    assign _1369 = !_1347;
    assign _1370 = _1369 & _1366;
    assign _1371 = _1368 | _1370;
    assign _1372 = _1332 | _1367;
    assign _1373 = _1332 & _1336;
    assign _1374 = !_1332;
    assign _1375 = _1374 & _1371;
    assign _1376 = _1373 | _1375;
    assign _1377 = _176 | _177;
    assign _1378 = _176 & _432;
    assign _1379 = !_176;
    assign _1380 = _1379 & _433;
    assign _1381 = _1378 | _1380;
    assign _1382 = _178 | _179;
    assign _1383 = _178 & _434;
    assign _1384 = !_178;
    assign _1385 = _1384 & _435;
    assign _1386 = _1383 | _1385;
    assign _1387 = _1377 | _1382;
    assign _1388 = _1377 & _1381;
    assign _1389 = !_1377;
    assign _1390 = _1389 & _1386;
    assign _1391 = _1388 | _1390;
    assign _1392 = _180 | _181;
    assign _1393 = _180 & _436;
    assign _1394 = !_180;
    assign _1395 = _1394 & _437;
    assign _1396 = _1393 | _1395;
    assign _1397 = _182 | _183;
    assign _1398 = _182 & _438;
    assign _1399 = !_182;
    assign _1400 = _1399 & _439;
    assign _1401 = _1398 | _1400;
    assign _1402 = _1392 | _1397;
    assign _1403 = _1392 & _1396;
    assign _1404 = !_1392;
    assign _1405 = _1404 & _1401;
    assign _1406 = _1403 | _1405;
    assign _1407 = _1387 | _1402;
    assign _1408 = _1387 & _1391;
    assign _1409 = !_1387;
    assign _1410 = _1409 & _1406;
    assign _1411 = _1408 | _1410;
    assign _1412 = _184 | _185;
    assign _1413 = _184 & _440;
    assign _1414 = !_184;
    assign _1415 = _1414 & _441;
    assign _1416 = _1413 | _1415;
    assign _1417 = _186 | _187;
    assign _1418 = _186 & _442;
    assign _1419 = !_186;
    assign _1420 = _1419 & _443;
    assign _1421 = _1418 | _1420;
    assign _1422 = _1412 | _1417;
    assign _1423 = _1412 & _1416;
    assign _1424 = !_1412;
    assign _1425 = _1424 & _1421;
    assign _1426 = _1423 | _1425;
    assign _1427 = _188 | _189;
    assign _1428 = _188 & _444;
    assign _1429 = !_188;
    assign _1430 = _1429 & _445;
    assign _1431 = _1428 | _1430;
    assign _1432 = _190 | _191;
    assign _1433 = _190 & _446;
    assign _1434 = !_190;
    assign _1435 = _1434 & _447;
    assign _1436 = _1433 | _1435;
    assign _1437 = _1427 | _1432;
    assign _1438 = _1427 & _1431;
    assign _1439 = !_1427;
    assign _1440 = _1439 & _1436;
    assign _1441 = _1438 | _1440;
    assign _1442 = _1422 | _1437;
    assign _1443 = _1422 & _1426;
    assign _1444 = !_1422;
    assign _1445 = _1444 & _1441;
    assign _1446 = _1443 | _1445;
    assign _1447 = _1407 | _1442;
    assign _1448 = _1407 & _1411;
    assign _1449 = !_1407;
    assign _1450 = _1449 & _1446;
    assign _1451 = _1448 | _1450;
    assign _1452 = _1372 | _1447;
    assign _1453 = _1372 & _1376;
    assign _1454 = !_1372;
    assign _1455 = _1454 & _1451;
    assign _1456 = _1453 | _1455;
    assign _1457 = _1297 | _1452;
    assign _1458 = _1297 & _1301;
    assign _1459 = !_1297;
    assign _1460 = _1459 & _1456;
    assign _1461 = _1458 | _1460;
    assign _1462 = _192 | _193;
    assign _1463 = _192 & _448;
    assign _1464 = !_192;
    assign _1465 = _1464 & _449;
    assign _1466 = _1463 | _1465;
    assign _1467 = _194 | _195;
    assign _1468 = _194 & _450;
    assign _1469 = !_194;
    assign _1470 = _1469 & _451;
    assign _1471 = _1468 | _1470;
    assign _1472 = _1462 | _1467;
    assign _1473 = _1462 & _1466;
    assign _1474 = !_1462;
    assign _1475 = _1474 & _1471;
    assign _1476 = _1473 | _1475;
    assign _1477 = _196 | _197;
    assign _1478 = _196 & _452;
    assign _1479 = !_196;
    assign _1480 = _1479 & _453;
    assign _1481 = _1478 | _1480;
    assign _1482 = _198 | _199;
    assign _1483 = _198 & _454;
    assign _1484 = !_198;
    assign _1485 = _1484 & _455;
    assign _1486 = _1483 | _1485;
    assign _1487 = _1477 | _1482;
    assign _1488 = _1477 & _1481;
    assign _1489 = !_1477;
    assign _1490 = _1489 & _1486;
    assign _1491 = _1488 | _1490;
    assign _1492 = _1472 | _1487;
    assign _1493 = _1472 & _1476;
    assign _1494 = !_1472;
    assign _1495 = _1494 & _1491;
    assign _1496 = _1493 | _1495;
    assign _1497 = _200 | _201;
    assign _1498 = _200 & _456;
    assign _1499 = !_200;
    assign _1500 = _1499 & _457;
    assign _1501 = _1498 | _1500;
    assign _1502 = _202 | _203;
    assign _1503 = _202 & _458;
    assign _1504 = !_202;
    assign _1505 = _1504 & _459;
    assign _1506 = _1503 | _1505;
    assign _1507 = _1497 | _1502;
    assign _1508 = _1497 & _1501;
    assign _1509 = !_1497;
    assign _1510 = _1509 & _1506;
    assign _1511 = _1508 | _1510;
    assign _1512 = _204 | _205;
    assign _1513 = _204 & _460;
    assign _1514 = !_204;
    assign _1515 = _1514 & _461;
    assign _1516 = _1513 | _1515;
    assign _1517 = _206 | _207;
    assign _1518 = _206 & _462;
    assign _1519 = !_206;
    assign _1520 = _1519 & _463;
    assign _1521 = _1518 | _1520;
    assign _1522 = _1512 | _1517;
    assign _1523 = _1512 & _1516;
    assign _1524 = !_1512;
    assign _1525 = _1524 & _1521;
    assign _1526 = _1523 | _1525;
    assign _1527 = _1507 | _1522;
    assign _1528 = _1507 & _1511;
    assign _1529 = !_1507;
    assign _1530 = _1529 & _1526;
    assign _1531 = _1528 | _1530;
    assign _1532 = _1492 | _1527;
    assign _1533 = _1492 & _1496;
    assign _1534 = !_1492;
    assign _1535 = _1534 & _1531;
    assign _1536 = _1533 | _1535;
    assign _1537 = _208 | _209;
    assign _1538 = _208 & _464;
    assign _1539 = !_208;
    assign _1540 = _1539 & _465;
    assign _1541 = _1538 | _1540;
    assign _1542 = _210 | _211;
    assign _1543 = _210 & _466;
    assign _1544 = !_210;
    assign _1545 = _1544 & _467;
    assign _1546 = _1543 | _1545;
    assign _1547 = _1537 | _1542;
    assign _1548 = _1537 & _1541;
    assign _1549 = !_1537;
    assign _1550 = _1549 & _1546;
    assign _1551 = _1548 | _1550;
    assign _1552 = _212 | _213;
    assign _1553 = _212 & _468;
    assign _1554 = !_212;
    assign _1555 = _1554 & _469;
    assign _1556 = _1553 | _1555;
    assign _1557 = _214 | _215;
    assign _1558 = _214 & _470;
    assign _1559 = !_214;
    assign _1560 = _1559 & _471;
    assign _1561 = _1558 | _1560;
    assign _1562 = _1552 | _1557;
    assign _1563 = _1552 & _1556;
    assign _1564 = !_1552;
    assign _1565 = _1564 & _1561;
    assign _1566 = _1563 | _1565;
    assign _1567 = _1547 | _1562;
    assign _1568 = _1547 & _1551;
    assign _1569 = !_1547;
    assign _1570 = _1569 & _1566;
    assign _1571 = _1568 | _1570;
    assign _1572 = _216 | _217;
    assign _1573 = _216 & _472;
    assign _1574 = !_216;
    assign _1575 = _1574 & _473;
    assign _1576 = _1573 | _1575;
    assign _1577 = _218 | _219;
    assign _1578 = _218 & _474;
    assign _1579 = !_218;
    assign _1580 = _1579 & _475;
    assign _1581 = _1578 | _1580;
    assign _1582 = _1572 | _1577;
    assign _1583 = _1572 & _1576;
    assign _1584 = !_1572;
    assign _1585 = _1584 & _1581;
    assign _1586 = _1583 | _1585;
    assign _1587 = _220 | _221;
    assign _1588 = _220 & _476;
    assign _1589 = !_220;
    assign _1590 = _1589 & _477;
    assign _1591 = _1588 | _1590;
    assign _1592 = _222 | _223;
    assign _1593 = _222 & _478;
    assign _1594 = !_222;
    assign _1595 = _1594 & _479;
    assign _1596 = _1593 | _1595;
    assign _1597 = _1587 | _1592;
    assign _1598 = _1587 & _1591;
    assign _1599 = !_1587;
    assign _1600 = _1599 & _1596;
    assign _1601 = _1598 | _1600;
    assign _1602 = _1582 | _1597;
    assign _1603 = _1582 & _1586;
    assign _1604 = !_1582;
    assign _1605 = _1604 & _1601;
    assign _1606 = _1603 | _1605;
    assign _1607 = _1567 | _1602;
    assign _1608 = _1567 & _1571;
    assign _1609 = !_1567;
    assign _1610 = _1609 & _1606;
    assign _1611 = _1608 | _1610;
    assign _1612 = _1532 | _1607;
    assign _1613 = _1532 & _1536;
    assign _1614 = !_1532;
    assign _1615 = _1614 & _1611;
    assign _1616 = _1613 | _1615;
    assign _1617 = _224 | _225;
    assign _1618 = _224 & _480;
    assign _1619 = !_224;
    assign _1620 = _1619 & _481;
    assign _1621 = _1618 | _1620;
    assign _1622 = _226 | _227;
    assign _1623 = _226 & _482;
    assign _1624 = !_226;
    assign _1625 = _1624 & _483;
    assign _1626 = _1623 | _1625;
    assign _1627 = _1617 | _1622;
    assign _1628 = _1617 & _1621;
    assign _1629 = !_1617;
    assign _1630 = _1629 & _1626;
    assign _1631 = _1628 | _1630;
    assign _1632 = _228 | _229;
    assign _1633 = _228 & _484;
    assign _1634 = !_228;
    assign _1635 = _1634 & _485;
    assign _1636 = _1633 | _1635;
    assign _1637 = _230 | _231;
    assign _1638 = _230 & _486;
    assign _1639 = !_230;
    assign _1640 = _1639 & _487;
    assign _1641 = _1638 | _1640;
    assign _1642 = _1632 | _1637;
    assign _1643 = _1632 & _1636;
    assign _1644 = !_1632;
    assign _1645 = _1644 & _1641;
    assign _1646 = _1643 | _1645;
    assign _1647 = _1627 | _1642;
    assign _1648 = _1627 & _1631;
    assign _1649 = !_1627;
    assign _1650 = _1649 & _1646;
    assign _1651 = _1648 | _1650;
    assign _1652 = _232 | _233;
    assign _1653 = _232 & _488;
    assign _1654 = !_232;
    assign _1655 = _1654 & _489;
    assign _1656 = _1653 | _1655;
    assign _1657 = _234 | _235;
    assign _1658 = _234 & _490;
    assign _1659 = !_234;
    assign _1660 = _1659 & _491;
    assign _1661 = _1658 | _1660;
    assign _1662 = _1652 | _1657;
    assign _1663 = _1652 & _1656;
    assign _1664 = !_1652;
    assign _1665 = _1664 & _1661;
    assign _1666 = _1663 | _1665;
    assign _1667 = _236 | _237;
    assign _1668 = _236 & _492;
    assign _1669 = !_236;
    assign _1670 = _1669 & _493;
    assign _1671 = _1668 | _1670;
    assign _1672 = _238 | _239;
    assign _1673 = _238 & _494;
    assign _1674 = !_238;
    assign _1675 = _1674 & _495;
    assign _1676 = _1673 | _1675;
    assign _1677 = _1667 | _1672;
    assign _1678 = _1667 & _1671;
    assign _1679 = !_1667;
    assign _1680 = _1679 & _1676;
    assign _1681 = _1678 | _1680;
    assign _1682 = _1662 | _1677;
    assign _1683 = _1662 & _1666;
    assign _1684 = !_1662;
    assign _1685 = _1684 & _1681;
    assign _1686 = _1683 | _1685;
    assign _1687 = _1647 | _1682;
    assign _1688 = _1647 & _1651;
    assign _1689 = !_1647;
    assign _1690 = _1689 & _1686;
    assign _1691 = _1688 | _1690;
    assign _1692 = _240 | _241;
    assign _1693 = _240 & _496;
    assign _1694 = !_240;
    assign _1695 = _1694 & _497;
    assign _1696 = _1693 | _1695;
    assign _1697 = _242 | _243;
    assign _1698 = _242 & _498;
    assign _1699 = !_242;
    assign _1700 = _1699 & _499;
    assign _1701 = _1698 | _1700;
    assign _1702 = _1692 | _1697;
    assign _1703 = _1692 & _1696;
    assign _1704 = !_1692;
    assign _1705 = _1704 & _1701;
    assign _1706 = _1703 | _1705;
    assign _1707 = _244 | _245;
    assign _1708 = _244 & _500;
    assign _1709 = !_244;
    assign _1710 = _1709 & _501;
    assign _1711 = _1708 | _1710;
    assign _1712 = _246 | _247;
    assign _1713 = _246 & _502;
    assign _1714 = !_246;
    assign _1715 = _1714 & _503;
    assign _1716 = _1713 | _1715;
    assign _1717 = _1707 | _1712;
    assign _1718 = _1707 & _1711;
    assign _1719 = !_1707;
    assign _1720 = _1719 & _1716;
    assign _1721 = _1718 | _1720;
    assign _1722 = _1702 | _1717;
    assign _1723 = _1702 & _1706;
    assign _1724 = !_1702;
    assign _1725 = _1724 & _1721;
    assign _1726 = _1723 | _1725;
    assign _1727 = _248 | _249;
    assign _1728 = _248 & _504;
    assign _1729 = !_248;
    assign _1730 = _1729 & _505;
    assign _1731 = _1728 | _1730;
    assign _1732 = _250 | _251;
    assign _1733 = _250 & _506;
    assign _1734 = !_250;
    assign _1735 = _1734 & _507;
    assign _1736 = _1733 | _1735;
    assign _1737 = _1727 | _1732;
    assign _1738 = _1727 & _1731;
    assign _1739 = !_1727;
    assign _1740 = _1739 & _1736;
    assign _1741 = _1738 | _1740;
    assign _1742 = _252 | _253;
    assign _1743 = _252 & _508;
    assign _1744 = !_252;
    assign _1745 = _1744 & _509;
    assign _1746 = _1743 | _1745;
    assign _1747 = _254 | _255;
    assign _1748 = _254 & _510;
    assign _1749 = !_254;
    assign _1750 = _1749 & _511;
    assign _1751 = _1748 | _1750;
    assign _1752 = _1742 | _1747;
    assign _1753 = _1742 & _1746;
    assign _1754 = !_1742;
    assign _1755 = _1754 & _1751;
    assign _1756 = _1753 | _1755;
    assign _1757 = _1737 | _1752;
    assign _1758 = _1737 & _1741;
    assign _1759 = !_1737;
    assign _1760 = _1759 & _1756;
    assign _1761 = _1758 | _1760;
    assign _1762 = _1722 | _1757;
    assign _1763 = _1722 & _1726;
    assign _1764 = !_1722;
    assign _1765 = _1764 & _1761;
    assign _1766 = _1763 | _1765;
    assign _1767 = _1687 | _1762;
    assign _1768 = _1687 & _1691;
    assign _1769 = !_1687;
    assign _1770 = _1769 & _1766;
    assign _1771 = _1768 | _1770;
    assign _1772 = _1612 | _1767;
    assign _1773 = _1612 & _1616;
    assign _1774 = !_1612;
    assign _1775 = _1774 & _1771;
    assign _1776 = _1773 | _1775;
    assign _1777 = _1457 | _1772;
    assign _1778 = _1457 & _1461;
    assign _1779 = !_1457;
    assign _1780 = _1779 & _1776;
    assign _1781 = _1778 | _1780;
    assign _1782 = _1142 | _1777;
    assign _1783 = _1142 & _1146;
    assign _1784 = !_1142;
    assign _1785 = _1784 & _1781;
    assign _1786 = _1783 | _1785;
    assign pp_ns = _1782;
    assign vv_ns = _1786;
    always @(posedge clk) begin
        pp <= pp_ns;
        vv <= vv_ns;
    end
endmodule

module swap(
    \a[0] ,
    \a[1] ,
    \a[2] ,
    \a[3] ,
    \a[4] ,
    \a[5] ,
    \a[6] ,
    \a[7] ,
    \a[8] ,
    \a[9] ,
    \a[10] ,
    \a[11] ,
    \a[12] ,
    \a[13] ,
    \a[14] ,
    \a[15] ,
    \b[0] ,
    \b[1] ,
    \b[2] ,
    \b[3] ,
    \b[4] ,
    \b[5] ,
    \b[6] ,
    \b[7] ,
    \b[8] ,
    \b[9] ,
    \b[10] ,
    \b[11] ,
    \b[12] ,
    \b[13] ,
    \b[14] ,
    \b[15] ,
    \x[0] ,
    \y[0] ,
    \x[1] ,
    \y[1] ,
    \x[2] ,
    \y[2] ,
    \x[3] ,
    \y[3] ,
    \x[4] ,
    \y[4] ,
    \x[5] ,
    \y[5] ,
    \x[6] ,
    \y[6] ,
    \x[7] ,
    \y[7] ,
    \x[8] ,
    \y[8] ,
    \x[9] ,
    \y[9] ,
    \x[10] ,
    \y[10] ,
    \x[11] ,
    \y[11] ,
    \x[12] ,
    \y[12] ,
    \x[13] ,
    \y[13] ,
    \x[14] ,
    \y[14] ,
    \x[15] ,
    \y[15] 
);
    input \a[0] ;
    input \a[1] ;
    input \a[2] ;
    input \a[3] ;
    input \a[4] ;
    input \a[5] ;
    input \a[6] ;
    input \a[7] ;
    input \a[8] ;
    input \a[9] ;
    input \a[10] ;
    input \a[11] ;
    input \a[12] ;
    input \a[13] ;
    input \a[14] ;
    input \a[15] ;
    input \b[0] ;
    input \b[1] ;
    input \b[2] ;
    input \b[3] ;
    input \b[4] ;
    input \b[5] ;
    input \b[6] ;
    input \b[7] ;
    input \b[8] ;
    input \b[9] ;
    input \b[10] ;
    input \b[11] ;
    input \b[12] ;
    input \b[13] ;
    input \b[14] ;
    input \b[15] ;
    output \x[0] ;
    output \y[0] ;
    output \x[1] ;
    output \y[1] ;
    output \x[2] ;
    output \y[2] ;
    output \x[3] ;
    output \y[3] ;
    output \x[4] ;
    output \y[4] ;
    output \x[5] ;
    output \y[5] ;
    output \x[6] ;
    output \y[6] ;
    output \x[7] ;
    output \y[7] ;
    output \x[8] ;
    output \y[8] ;
    output \x[9] ;
    output \y[9] ;
    output \x[10] ;
    output \y[10] ;
    output \x[11] ;
    output \y[11] ;
    output \x[12] ;
    output \y[12] ;
    output \x[13] ;
    output \y[13] ;
    output \x[14] ;
    output \y[14] ;
    output \x[15] ;
    output \y[15] ;
    wire _0;
    wire _1;
    wire _2;
    wire _3;
    wire _4;
    wire _5;
    wire _6;
    wire _7;
    wire _8;
    wire _9;
    wire _10;
    wire _11;
    wire _12;
    wire _13;
    wire _14;
    wire _15;
    wire _16;
    wire _17;
    wire _18;
    wire _19;
    wire _20;
    wire _21;
    wire _22;
    wire _23;
    wire _24;
    wire _25;
    wire _26;
    wire _27;
    wire _28;
    wire _29;
    wire _30;
    wire _31;
    wire _32;
    wire _33;
    wire _34;
    wire _35;
    wire _36;
    wire _37;
    wire _38;
    wire _39;
    wire _40;
    wire _41;
    wire _42;
    wire _43;
    wire _44;
    wire _45;
    wire _46;
    wire _47;
    wire _48;
    wire _49;
    wire _50;
    wire _51;
    wire _52;
    wire _53;
    wire _54;
    wire _55;
    wire _56;
    wire _57;
    wire _58;
    wire _59;
    wire _60;
    wire _61;
    wire _62;
    wire _63;
    wire _64;
    wire _65;
    wire _66;
    wire _67;
    wire _68;
    wire _69;
    wire _70;
    wire _71;
    wire _72;
    wire _73;
    wire _74;
    wire _75;
    wire _76;
    wire _77;
    wire _78;
    wire _79;
    wire _80;
    wire _81;
    wire _82;
    wire _83;
    wire _84;
    wire _85;
    wire _86;
    wire _87;
    wire _88;
    wire _89;
    wire _90;
    wire _91;
    wire _92;
    wire _93;
    wire _94;
    wire _95;
    wire _96;
    wire _97;
    wire _98;
    wire _99;
    wire _100;
    wire _101;
    wire _102;
    wire _103;
    wire _104;
    wire _105;
    wire _106;
    wire _107;
    wire _108;
    wire _109;
    wire _110;
    wire _111;
    wire _112;
    wire _113;
    wire _114;
    wire _115;
    wire _116;
    wire _117;
    wire _118;
    wire _119;
    wire _120;
    wire _121;
    wire _122;
    wire _123;
    wire _124;
    wire _125;
    wire _126;
    wire _127;
    wire _128;
    wire _129;
    wire _130;
    wire _131;
    wire _132;
    wire _133;
    wire _134;
    wire _135;
    wire _136;
    wire _137;
    wire _138;
    wire _139;
    wire _140;
    wire _141;
    wire _142;
    wire _143;
    wire _144;
    wire _145;
    wire _146;
    wire _147;
    wire _148;
    wire _149;
    wire _150;
    wire _151;
    wire _152;
    wire _153;
    wire _154;
    wire _155;
    wire _156;
    wire _157;
    wire _158;
    wire _159;
    wire _160;
    wire _161;
    wire _162;
    wire _163;
    wire _164;
    wire _165;
    wire _166;
    wire _167;
    wire _168;
    wire _169;
    wire _170;
    wire _171;
    wire _172;
    wire _173;
    wire _174;
    wire _175;
    wire _176;
    wire _177;
    wire _178;
    wire _179;
    wire _180;
    wire _181;
    wire _182;
    wire _183;
    wire _184;
    wire _185;
    wire _186;
    wire _187;
    wire _188;
    wire _189;
    wire _190;
    wire _191;
    wire _192;
    wire _193;
    wire _194;
    wire _195;
    wire _196;
    wire _197;
    wire _198;
    wire _199;
    wire _200;
    wire _201;
    wire _202;
    wire _203;
    wire _204;
    wire _205;
    wire _206;
    wire _207;
    wire _208;
    wire _209;
    wire _210;
    wire _211;
    wire _212;
    wire _213;
    wire _214;
    wire _215;
    wire _216;
    wire _217;
    wire _218;
    wire _219;
    wire _220;
    wire _221;
    wire _222;
    wire _223;
    wire _224;
    wire _225;
    wire _226;
    wire _227;
    wire _228;
    wire _229;
    wire _230;
    wire _231;
    wire _232;
    wire _233;
    wire _234;
    wire _235;
    wire _236;
    wire _237;
    wire _238;
    wire _239;
    wire _240;
    wire _241;
    wire _242;
    wire _243;
    wire _244;
    wire _245;
    wire _246;
    wire _247;
    wire _248;
    wire _249;
    wire _250;
    wire _251;
    wire _252;
    wire _253;
    wire _254;
    wire _255;
    wire _256;
    wire _257;
    wire _258;
    wire _259;
    wire _260;
    wire _261;
    wire _262;
    wire _263;
    wire _264;
    wire _265;
    wire _266;
    wire _267;
    wire _268;
    wire _269;
    wire _270;
    wire _271;
    wire _272;
    wire _273;
    wire _274;
    wire _275;
    wire _276;
    wire _277;
    wire _278;
    wire _279;
    wire _280;
    wire _281;
    wire _282;
    wire _283;
    wire _284;
    wire _285;
    wire _286;
    wire _287;
    wire _288;
    wire _289;
    wire _290;
    wire _291;
    wire _292;
    wire _293;
    wire _294;
    wire _295;
    wire _296;
    wire _297;
    wire _298;
    wire _299;
    wire _300;
    wire _301;
    wire _302;
    wire _303;
    wire _304;
    wire _305;
    wire _306;
    wire _307;
    wire _308;
    wire _309;
    wire _310;
    wire _311;
    wire _312;
    wire _313;
    wire _314;
    wire _315;
    wire _316;
    wire _317;
    assign _0 = \a[0] ;
    assign _1 = \a[1] ;
    assign _2 = \a[2] ;
    assign _3 = \a[3] ;
    assign _4 = \a[4] ;
    assign _5 = \a[5] ;
    assign _6 = \a[6] ;
    assign _7 = \a[7] ;
    assign _8 = \a[8] ;
    assign _9 = \a[9] ;
    assign _10 = \a[10] ;
    assign _11 = \a[11] ;
    assign _12 = \a[12] ;
    assign _13 = \a[13] ;
    assign _14 = \a[14] ;
    assign _15 = \a[15] ;
    assign _16 = \b[0] ;
    assign _17 = \b[1] ;
    assign _18 = \b[2] ;
    assign _19 = \b[3] ;
    assign _20 = \b[4] ;
    assign _21 = \b[5] ;
    assign _22 = \b[6] ;
    assign _23 = \b[7] ;
    assign _24 = \b[8] ;
    assign _25 = \b[9] ;
    assign _26 = \b[10] ;
    assign _27 = \b[11] ;
    assign _28 = \b[12] ;
    assign _29 = \b[13] ;
    assign _30 = \b[14] ;
    assign _31 = \b[15] ;
    assign _32 = !_0;
    assign _33 = _32 & _16;
    assign _34 = !_0;
    assign _35 = !_16;
    assign _36 = _34 & _35;
    assign _37 = _0 & _16;
    assign _38 = _36 | _37;
    assign _39 = !_1;
    assign _40 = _39 & _17;
    assign _41 = !_1;
    assign _42 = !_17;
    assign _43 = _41 & _42;
    assign _44 = _1 & _17;
    assign _45 = _43 | _44;
    assign _46 = _45 & _33;
    assign _47 = _40 | _46;
    assign _48 = _45 & _38;
    assign _49 = !_2;
    assign _50 = _49 & _18;
    assign _51 = !_2;
    assign _52 = !_18;
    assign _53 = _51 & _52;
    assign _54 = _2 & _18;
    assign _55 = _53 | _54;
    assign _56 = !_3;
    assign _57 = _56 & _19;
    assign _58 = !_3;
    assign _59 = !_19;
    assign _60 = _58 & _59;
    assign _61 = _3 & _19;
    assign _62 = _60 | _61;
    assign _63 = _62 & _50;
    assign _64 = _57 | _63;
    assign _65 = _62 & _55;
    assign _66 = _65 & _47;
    assign _67 = _64 | _66;
    assign _68 = _65 & _48;
    assign _69 = !_4;
    assign _70 = _69 & _20;
    assign _71 = !_4;
    assign _72 = !_20;
    assign _73 = _71 & _72;
    assign _74 = _4 & _20;
    assign _75 = _73 | _74;
    assign _76 = !_5;
    assign _77 = _76 & _21;
    assign _78 = !_5;
    assign _79 = !_21;
    assign _80 = _78 & _79;
    assign _81 = _5 & _21;
    assign _82 = _80 | _81;
    assign _83 = _82 & _70;
    assign _84 = _77 | _83;
    assign _85 = _82 & _75;
    assign _86 = !_6;
    assign _87 = _86 & _22;
    assign _88 = !_6;
    assign _89 = !_22;
    assign _90 = _88 & _89;
    assign _91 = _6 & _22;
    assign _92 = _90 | _91;
    assign _93 = !_7;
    assign _94 = _93 & _23;
    assign _95 = !_7;
    assign _96 = !_23;
    assign _97 = _95 & _96;
    assign _98 = _7 & _23;
    assign _99 = _97 | _98;
    assign _100 = _99 & _87;
    assign _101 = _94 | _100;
    assign _102 = _99 & _92;
    assign _103 = _102 & _84;
    assign _104 = _101 | _103;
    assign _105 = _102 & _85;
    assign _106 = _105 & _67;
    assign _107 = _104 | _106;
    assign _108 = _105 & _68;
    assign _109 = !_8;
    assign _110 = _109 & _24;
    assign _111 = !_8;
    assign _112 = !_24;
    assign _113 = _111 & _112;
    assign _114 = _8 & _24;
    assign _115 = _113 | _114;
    assign _116 = !_9;
    assign _117 = _116 & _25;
    assign _118 = !_9;
    assign _119 = !_25;
    assign _120 = _118 & _119;
    assign _121 = _9 & _25;
    assign _122 = _120 | _121;
    assign _123 = _122 & _110;
    assign _124 = _117 | _123;
    assign _125 = _122 & _115;
    assign _126 = !_10;
    assign _127 = _126 & _26;
    assign _128 = !_10;
    assign _129 = !_26;
    assign _130 = _128 & _129;
    assign _131 = _10 & _26;
    assign _132 = _130 | _131;
    assign _133 = !_11;
    assign _134 = _133 & _27;
    assign _135 = !_11;
    assign _136 = !_27;
    assign _137 = _135 & _136;
    assign _138 = _11 & _27;
    assign _139 = _137 | _138;
    assign _140 = _139 & _127;
    assign _141 = _134 | _140;
    assign _142 = _139 & _132;
    assign _143 = _142 & _124;
    assign _144 = _141 | _143;
    assign _145 = _142 & _125;
    assign _146 = !_12;
    assign _147 = _146 & _28;
    assign _148 = !_12;
    assign _149 = !_28;
    assign _150 = _148 & _149;
    assign _151 = _12 & _28;
    assign _152 = _150 | _151;
    assign _153 = !_13;
    assign _154 = _153 & _29;
    assign _155 = !_13;
    assign _156 = !_29;
    assign _157 = _155 & _156;
    assign _158 = _13 & _29;
    assign _159 = _157 | _158;
    assign _160 = _159 & _147;
    assign _161 = _154 | _160;
    assign _162 = _159 & _152;
    assign _163 = !_14;
    assign _164 = _163 & _30;
    assign _165 = !_14;
    assign _166 = !_30;
    assign _167 = _165 & _166;
    assign _168 = _14 & _30;
    assign _169 = _167 | _168;
    assign _170 = !_15;
    assign _171 = _170 & _31;
    assign _172 = !_15;
    assign _173 = !_31;
    assign _174 = _172 & _173;
    assign _175 = _15 & _31;
    assign _176 = _174 | _175;
    assign _177 = _176 & _164;
    assign _178 = _171 | _177;
    assign _179 = _176 & _169;
    assign _180 = _179 & _161;
    assign _181 = _178 | _180;
    assign _182 = _179 & _162;
    assign _183 = _182 & _144;
    assign _184 = _181 | _183;
    assign _185 = _182 & _145;
    assign _186 = _185 & _107;
    assign _187 = _184 | _186;
    assign _188 = _185 & _108;
    assign _189 = _187 & _0;
    assign _190 = !_187;
    assign _191 = _190 & _16;
    assign _192 = _189 | _191;
    assign _193 = _187 & _1;
    assign _194 = !_187;
    assign _195 = _194 & _17;
    assign _196 = _193 | _195;
    assign _197 = _187 & _2;
    assign _198 = !_187;
    assign _199 = _198 & _18;
    assign _200 = _197 | _199;
    assign _201 = _187 & _3;
    assign _202 = !_187;
    assign _203 = _202 & _19;
    assign _204 = _201 | _203;
    assign _205 = _187 & _4;
    assign _206 = !_187;
    assign _207 = _206 & _20;
    assign _208 = _205 | _207;
    assign _209 = _187 & _5;
    assign _210 = !_187;
    assign _211 = _210 & _21;
    assign _212 = _209 | _211;
    assign _213 = _187 & _6;
    assign _214 = !_187;
    assign _215 = _214 & _22;
    assign _216 = _213 | _215;
    assign _217 = _187 & _7;
    assign _218 = !_187;
    assign _219 = _218 & _23;
    assign _220 = _217 | _219;
    assign _221 = _187 & _8;
    assign _222 = !_187;
    assign _223 = _222 & _24;
    assign _224 = _221 | _223;
    assign _225 = _187 & _9;
    assign _226 = !_187;
    assign _227 = _226 & _25;
    assign _228 = _225 | _227;
    assign _229 = _187 & _10;
    assign _230 = !_187;
    assign _231 = _230 & _26;
    assign _232 = _229 | _231;
    assign _233 = _187 & _11;
    assign _234 = !_187;
    assign _235 = _234 & _27;
    assign _236 = _233 | _235;
    assign _237 = _187 & _12;
    assign _238 = !_187;
    assign _239 = _238 & _28;
    assign _240 = _237 | _239;
    assign _241 = _187 & _13;
    assign _242 = !_187;
    assign _243 = _242 & _29;
    assign _244 = _241 | _243;
    assign _245 = _187 & _14;
    assign _246 = !_187;
    assign _247 = _246 & _30;
    assign _248 = _245 | _247;
    assign _249 = _187 & _15;
    assign _250 = !_187;
    assign _251 = _250 & _31;
    assign _252 = _249 | _251;
    assign _253 = !_187;
    assign _254 = _253 & _0;
    assign _255 = !_253;
    assign _256 = _255 & _16;
    assign _257 = _254 | _256;
    assign _258 = _253 & _1;
    assign _259 = !_253;
    assign _260 = _259 & _17;
    assign _261 = _258 | _260;
    assign _262 = _253 & _2;
    assign _263 = !_253;
    assign _264 = _263 & _18;
    assign _265 = _262 | _264;
    assign _266 = _253 & _3;
    assign _267 = !_253;
    assign _268 = _267 & _19;
    assign _269 = _266 | _268;
    assign _270 = _253 & _4;
    assign _271 = !_253;
    assign _272 = _271 & _20;
    assign _273 = _270 | _272;
    assign _274 = _253 & _5;
    assign _275 = !_253;
    assign _276 = _275 & _21;
    assign _277 = _274 | _276;
    assign _278 = _253 & _6;
    assign _279 = !_253;
    assign _280 = _279 & _22;
    assign _281 = _278 | _280;
    assign _282 = _253 & _7;
    assign _283 = !_253;
    assign _284 = _283 & _23;
    assign _285 = _282 | _284;
    assign _286 = _253 & _8;
    assign _287 = !_253;
    assign _288 = _287 & _24;
    assign _289 = _286 | _288;
    assign _290 = _253 & _9;
    assign _291 = !_253;
    assign _292 = _291 & _25;
    assign _293 = _290 | _292;
    assign _294 = _253 & _10;
    assign _295 = !_253;
    assign _296 = _295 & _26;
    assign _297 = _294 | _296;
    assign _298 = _253 & _11;
    assign _299 = !_253;
    assign _300 = _299 & _27;
    assign _301 = _298 | _300;
    assign _302 = _253 & _12;
    assign _303 = !_253;
    assign _304 = _303 & _28;
    assign _305 = _302 | _304;
    assign _306 = _253 & _13;
    assign _307 = !_253;
    assign _308 = _307 & _29;
    assign _309 = _306 | _308;
    assign _310 = _253 & _14;
    assign _311 = !_253;
    assign _312 = _311 & _30;
    assign _313 = _310 | _312;
    assign _314 = _253 & _15;
    assign _315 = !_253;
    assign _316 = _315 & _31;
    assign _317 = _314 | _316;
    assign \x[0]  = _192;
    assign \y[0]  = _257;
    assign \x[1]  = _196;
    assign \y[1]  = _261;
    assign \x[2]  = _200;
    assign \y[2]  = _265;
    assign \x[3]  = _204;
    assign \y[3]  = _269;
    assign \x[4]  = _208;
    assign \y[4]  = _273;
    assign \x[5]  = _212;
    assign \y[5]  = _277;
    assign \x[6]  = _216;
    assign \y[6]  = _281;
    assign \x[7]  = _220;
    assign \y[7]  = _285;
    assign \x[8]  = _224;
    assign \y[8]  = _289;
    assign \x[9]  = _228;
    assign \y[9]  = _293;
    assign \x[10]  = _232;
    assign \y[10]  = _297;
    assign \x[11]  = _236;
    assign \y[11]  = _301;
    assign \x[12]  = _240;
    assign \y[12]  = _305;
    assign \x[13]  = _244;
    assign \y[13]  = _309;
    assign \x[14]  = _248;
    assign \y[14]  = _313;
    assign \x[15]  = _252;
    assign \y[15]  = _317;
endmodule

module bitonic_recursive(
    \a[0][0] ,
    \a[0][1] ,
    \a[0][2] ,
    \a[0][3] ,
    \a[0][4] ,
    \a[0][5] ,
    \a[0][6] ,
    \a[0][7] ,
    \a[0][8] ,
    \a[0][9] ,
    \a[0][10] ,
    \a[0][11] ,
    \a[0][12] ,
    \a[0][13] ,
    \a[0][14] ,
    \a[0][15] ,
    \a[1][0] ,
    \a[1][1] ,
    \a[1][2] ,
    \a[1][3] ,
    \a[1][4] ,
    \a[1][5] ,
    \a[1][6] ,
    \a[1][7] ,
    \a[1][8] ,
    \a[1][9] ,
    \a[1][10] ,
    \a[1][11] ,
    \a[1][12] ,
    \a[1][13] ,
    \a[1][14] ,
    \a[1][15] ,
    \a[2][0] ,
    \a[2][1] ,
    \a[2][2] ,
    \a[2][3] ,
    \a[2][4] ,
    \a[2][5] ,
    \a[2][6] ,
    \a[2][7] ,
    \a[2][8] ,
    \a[2][9] ,
    \a[2][10] ,
    \a[2][11] ,
    \a[2][12] ,
    \a[2][13] ,
    \a[2][14] ,
    \a[2][15] ,
    \a[3][0] ,
    \a[3][1] ,
    \a[3][2] ,
    \a[3][3] ,
    \a[3][4] ,
    \a[3][5] ,
    \a[3][6] ,
    \a[3][7] ,
    \a[3][8] ,
    \a[3][9] ,
    \a[3][10] ,
    \a[3][11] ,
    \a[3][12] ,
    \a[3][13] ,
    \a[3][14] ,
    \a[3][15] ,
    \a[4][0] ,
    \a[4][1] ,
    \a[4][2] ,
    \a[4][3] ,
    \a[4][4] ,
    \a[4][5] ,
    \a[4][6] ,
    \a[4][7] ,
    \a[4][8] ,
    \a[4][9] ,
    \a[4][10] ,
    \a[4][11] ,
    \a[4][12] ,
    \a[4][13] ,
    \a[4][14] ,
    \a[4][15] ,
    \a[5][0] ,
    \a[5][1] ,
    \a[5][2] ,
    \a[5][3] ,
    \a[5][4] ,
    \a[5][5] ,
    \a[5][6] ,
    \a[5][7] ,
    \a[5][8] ,
    \a[5][9] ,
    \a[5][10] ,
    \a[5][11] ,
    \a[5][12] ,
    \a[5][13] ,
    \a[5][14] ,
    \a[5][15] ,
    \a[6][0] ,
    \a[6][1] ,
    \a[6][2] ,
    \a[6][3] ,
    \a[6][4] ,
    \a[6][5] ,
    \a[6][6] ,
    \a[6][7] ,
    \a[6][8] ,
    \a[6][9] ,
    \a[6][10] ,
    \a[6][11] ,
    \a[6][12] ,
    \a[6][13] ,
    \a[6][14] ,
    \a[6][15] ,
    \a[7][0] ,
    \a[7][1] ,
    \a[7][2] ,
    \a[7][3] ,
    \a[7][4] ,
    \a[7][5] ,
    \a[7][6] ,
    \a[7][7] ,
    \a[7][8] ,
    \a[7][9] ,
    \a[7][10] ,
    \a[7][11] ,
    \a[7][12] ,
    \a[7][13] ,
    \a[7][14] ,
    \a[7][15] ,
    \a[8][0] ,
    \a[8][1] ,
    \a[8][2] ,
    \a[8][3] ,
    \a[8][4] ,
    \a[8][5] ,
    \a[8][6] ,
    \a[8][7] ,
    \a[8][8] ,
    \a[8][9] ,
    \a[8][10] ,
    \a[8][11] ,
    \a[8][12] ,
    \a[8][13] ,
    \a[8][14] ,
    \a[8][15] ,
    \a[9][0] ,
    \a[9][1] ,
    \a[9][2] ,
    \a[9][3] ,
    \a[9][4] ,
    \a[9][5] ,
    \a[9][6] ,
    \a[9][7] ,
    \a[9][8] ,
    \a[9][9] ,
    \a[9][10] ,
    \a[9][11] ,
    \a[9][12] ,
    \a[9][13] ,
    \a[9][14] ,
    \a[9][15] ,
    \a[10][0] ,
    \a[10][1] ,
    \a[10][2] ,
    \a[10][3] ,
    \a[10][4] ,
    \a[10][5] ,
    \a[10][6] ,
    \a[10][7] ,
    \a[10][8] ,
    \a[10][9] ,
    \a[10][10] ,
    \a[10][11] ,
    \a[10][12] ,
    \a[10][13] ,
    \a[10][14] ,
    \a[10][15] ,
    \a[11][0] ,
    \a[11][1] ,
    \a[11][2] ,
    \a[11][3] ,
    \a[11][4] ,
    \a[11][5] ,
    \a[11][6] ,
    \a[11][7] ,
    \a[11][8] ,
    \a[11][9] ,
    \a[11][10] ,
    \a[11][11] ,
    \a[11][12] ,
    \a[11][13] ,
    \a[11][14] ,
    \a[11][15] ,
    \a[12][0] ,
    \a[12][1] ,
    \a[12][2] ,
    \a[12][3] ,
    \a[12][4] ,
    \a[12][5] ,
    \a[12][6] ,
    \a[12][7] ,
    \a[12][8] ,
    \a[12][9] ,
    \a[12][10] ,
    \a[12][11] ,
    \a[12][12] ,
    \a[12][13] ,
    \a[12][14] ,
    \a[12][15] ,
    \a[13][0] ,
    \a[13][1] ,
    \a[13][2] ,
    \a[13][3] ,
    \a[13][4] ,
    \a[13][5] ,
    \a[13][6] ,
    \a[13][7] ,
    \a[13][8] ,
    \a[13][9] ,
    \a[13][10] ,
    \a[13][11] ,
    \a[13][12] ,
    \a[13][13] ,
    \a[13][14] ,
    \a[13][15] ,
    \a[14][0] ,
    \a[14][1] ,
    \a[14][2] ,
    \a[14][3] ,
    \a[14][4] ,
    \a[14][5] ,
    \a[14][6] ,
    \a[14][7] ,
    \a[14][8] ,
    \a[14][9] ,
    \a[14][10] ,
    \a[14][11] ,
    \a[14][12] ,
    \a[14][13] ,
    \a[14][14] ,
    \a[14][15] ,
    \a[15][0] ,
    \a[15][1] ,
    \a[15][2] ,
    \a[15][3] ,
    \a[15][4] ,
    \a[15][5] ,
    \a[15][6] ,
    \a[15][7] ,
    \a[15][8] ,
    \a[15][9] ,
    \a[15][10] ,
    \a[15][11] ,
    \a[15][12] ,
    \a[15][13] ,
    \a[15][14] ,
    \a[15][15] ,
    \a_sorted[0][0] ,
    \a_sorted[0][1] ,
    \a_sorted[0][2] ,
    \a_sorted[0][3] ,
    \a_sorted[0][4] ,
    \a_sorted[0][5] ,
    \a_sorted[0][6] ,
    \a_sorted[0][7] ,
    \a_sorted[0][8] ,
    \a_sorted[0][9] ,
    \a_sorted[0][10] ,
    \a_sorted[0][11] ,
    \a_sorted[0][12] ,
    \a_sorted[0][13] ,
    \a_sorted[0][14] ,
    \a_sorted[0][15] ,
    \a_sorted[1][0] ,
    \a_sorted[1][1] ,
    \a_sorted[1][2] ,
    \a_sorted[1][3] ,
    \a_sorted[1][4] ,
    \a_sorted[1][5] ,
    \a_sorted[1][6] ,
    \a_sorted[1][7] ,
    \a_sorted[1][8] ,
    \a_sorted[1][9] ,
    \a_sorted[1][10] ,
    \a_sorted[1][11] ,
    \a_sorted[1][12] ,
    \a_sorted[1][13] ,
    \a_sorted[1][14] ,
    \a_sorted[1][15] ,
    \a_sorted[2][0] ,
    \a_sorted[2][1] ,
    \a_sorted[2][2] ,
    \a_sorted[2][3] ,
    \a_sorted[2][4] ,
    \a_sorted[2][5] ,
    \a_sorted[2][6] ,
    \a_sorted[2][7] ,
    \a_sorted[2][8] ,
    \a_sorted[2][9] ,
    \a_sorted[2][10] ,
    \a_sorted[2][11] ,
    \a_sorted[2][12] ,
    \a_sorted[2][13] ,
    \a_sorted[2][14] ,
    \a_sorted[2][15] ,
    \a_sorted[3][0] ,
    \a_sorted[3][1] ,
    \a_sorted[3][2] ,
    \a_sorted[3][3] ,
    \a_sorted[3][4] ,
    \a_sorted[3][5] ,
    \a_sorted[3][6] ,
    \a_sorted[3][7] ,
    \a_sorted[3][8] ,
    \a_sorted[3][9] ,
    \a_sorted[3][10] ,
    \a_sorted[3][11] ,
    \a_sorted[3][12] ,
    \a_sorted[3][13] ,
    \a_sorted[3][14] ,
    \a_sorted[3][15] ,
    \a_sorted[4][0] ,
    \a_sorted[4][1] ,
    \a_sorted[4][2] ,
    \a_sorted[4][3] ,
    \a_sorted[4][4] ,
    \a_sorted[4][5] ,
    \a_sorted[4][6] ,
    \a_sorted[4][7] ,
    \a_sorted[4][8] ,
    \a_sorted[4][9] ,
    \a_sorted[4][10] ,
    \a_sorted[4][11] ,
    \a_sorted[4][12] ,
    \a_sorted[4][13] ,
    \a_sorted[4][14] ,
    \a_sorted[4][15] ,
    \a_sorted[5][0] ,
    \a_sorted[5][1] ,
    \a_sorted[5][2] ,
    \a_sorted[5][3] ,
    \a_sorted[5][4] ,
    \a_sorted[5][5] ,
    \a_sorted[5][6] ,
    \a_sorted[5][7] ,
    \a_sorted[5][8] ,
    \a_sorted[5][9] ,
    \a_sorted[5][10] ,
    \a_sorted[5][11] ,
    \a_sorted[5][12] ,
    \a_sorted[5][13] ,
    \a_sorted[5][14] ,
    \a_sorted[5][15] ,
    \a_sorted[6][0] ,
    \a_sorted[6][1] ,
    \a_sorted[6][2] ,
    \a_sorted[6][3] ,
    \a_sorted[6][4] ,
    \a_sorted[6][5] ,
    \a_sorted[6][6] ,
    \a_sorted[6][7] ,
    \a_sorted[6][8] ,
    \a_sorted[6][9] ,
    \a_sorted[6][10] ,
    \a_sorted[6][11] ,
    \a_sorted[6][12] ,
    \a_sorted[6][13] ,
    \a_sorted[6][14] ,
    \a_sorted[6][15] ,
    \a_sorted[7][0] ,
    \a_sorted[7][1] ,
    \a_sorted[7][2] ,
    \a_sorted[7][3] ,
    \a_sorted[7][4] ,
    \a_sorted[7][5] ,
    \a_sorted[7][6] ,
    \a_sorted[7][7] ,
    \a_sorted[7][8] ,
    \a_sorted[7][9] ,
    \a_sorted[7][10] ,
    \a_sorted[7][11] ,
    \a_sorted[7][12] ,
    \a_sorted[7][13] ,
    \a_sorted[7][14] ,
    \a_sorted[7][15] ,
    \a_sorted[8][0] ,
    \a_sorted[8][1] ,
    \a_sorted[8][2] ,
    \a_sorted[8][3] ,
    \a_sorted[8][4] ,
    \a_sorted[8][5] ,
    \a_sorted[8][6] ,
    \a_sorted[8][7] ,
    \a_sorted[8][8] ,
    \a_sorted[8][9] ,
    \a_sorted[8][10] ,
    \a_sorted[8][11] ,
    \a_sorted[8][12] ,
    \a_sorted[8][13] ,
    \a_sorted[8][14] ,
    \a_sorted[8][15] ,
    \a_sorted[9][0] ,
    \a_sorted[9][1] ,
    \a_sorted[9][2] ,
    \a_sorted[9][3] ,
    \a_sorted[9][4] ,
    \a_sorted[9][5] ,
    \a_sorted[9][6] ,
    \a_sorted[9][7] ,
    \a_sorted[9][8] ,
    \a_sorted[9][9] ,
    \a_sorted[9][10] ,
    \a_sorted[9][11] ,
    \a_sorted[9][12] ,
    \a_sorted[9][13] ,
    \a_sorted[9][14] ,
    \a_sorted[9][15] ,
    \a_sorted[10][0] ,
    \a_sorted[10][1] ,
    \a_sorted[10][2] ,
    \a_sorted[10][3] ,
    \a_sorted[10][4] ,
    \a_sorted[10][5] ,
    \a_sorted[10][6] ,
    \a_sorted[10][7] ,
    \a_sorted[10][8] ,
    \a_sorted[10][9] ,
    \a_sorted[10][10] ,
    \a_sorted[10][11] ,
    \a_sorted[10][12] ,
    \a_sorted[10][13] ,
    \a_sorted[10][14] ,
    \a_sorted[10][15] ,
    \a_sorted[11][0] ,
    \a_sorted[11][1] ,
    \a_sorted[11][2] ,
    \a_sorted[11][3] ,
    \a_sorted[11][4] ,
    \a_sorted[11][5] ,
    \a_sorted[11][6] ,
    \a_sorted[11][7] ,
    \a_sorted[11][8] ,
    \a_sorted[11][9] ,
    \a_sorted[11][10] ,
    \a_sorted[11][11] ,
    \a_sorted[11][12] ,
    \a_sorted[11][13] ,
    \a_sorted[11][14] ,
    \a_sorted[11][15] ,
    \a_sorted[12][0] ,
    \a_sorted[12][1] ,
    \a_sorted[12][2] ,
    \a_sorted[12][3] ,
    \a_sorted[12][4] ,
    \a_sorted[12][5] ,
    \a_sorted[12][6] ,
    \a_sorted[12][7] ,
    \a_sorted[12][8] ,
    \a_sorted[12][9] ,
    \a_sorted[12][10] ,
    \a_sorted[12][11] ,
    \a_sorted[12][12] ,
    \a_sorted[12][13] ,
    \a_sorted[12][14] ,
    \a_sorted[12][15] ,
    \a_sorted[13][0] ,
    \a_sorted[13][1] ,
    \a_sorted[13][2] ,
    \a_sorted[13][3] ,
    \a_sorted[13][4] ,
    \a_sorted[13][5] ,
    \a_sorted[13][6] ,
    \a_sorted[13][7] ,
    \a_sorted[13][8] ,
    \a_sorted[13][9] ,
    \a_sorted[13][10] ,
    \a_sorted[13][11] ,
    \a_sorted[13][12] ,
    \a_sorted[13][13] ,
    \a_sorted[13][14] ,
    \a_sorted[13][15] ,
    \a_sorted[14][0] ,
    \a_sorted[14][1] ,
    \a_sorted[14][2] ,
    \a_sorted[14][3] ,
    \a_sorted[14][4] ,
    \a_sorted[14][5] ,
    \a_sorted[14][6] ,
    \a_sorted[14][7] ,
    \a_sorted[14][8] ,
    \a_sorted[14][9] ,
    \a_sorted[14][10] ,
    \a_sorted[14][11] ,
    \a_sorted[14][12] ,
    \a_sorted[14][13] ,
    \a_sorted[14][14] ,
    \a_sorted[14][15] ,
    \a_sorted[15][0] ,
    \a_sorted[15][1] ,
    \a_sorted[15][2] ,
    \a_sorted[15][3] ,
    \a_sorted[15][4] ,
    \a_sorted[15][5] ,
    \a_sorted[15][6] ,
    \a_sorted[15][7] ,
    \a_sorted[15][8] ,
    \a_sorted[15][9] ,
    \a_sorted[15][10] ,
    \a_sorted[15][11] ,
    \a_sorted[15][12] ,
    \a_sorted[15][13] ,
    \a_sorted[15][14] ,
    \a_sorted[15][15] ,
    clk
);
    input clk;
    input \a[0][0] ;
    input \a[0][1] ;
    input \a[0][2] ;
    input \a[0][3] ;
    input \a[0][4] ;
    input \a[0][5] ;
    input \a[0][6] ;
    input \a[0][7] ;
    input \a[0][8] ;
    input \a[0][9] ;
    input \a[0][10] ;
    input \a[0][11] ;
    input \a[0][12] ;
    input \a[0][13] ;
    input \a[0][14] ;
    input \a[0][15] ;
    input \a[1][0] ;
    input \a[1][1] ;
    input \a[1][2] ;
    input \a[1][3] ;
    input \a[1][4] ;
    input \a[1][5] ;
    input \a[1][6] ;
    input \a[1][7] ;
    input \a[1][8] ;
    input \a[1][9] ;
    input \a[1][10] ;
    input \a[1][11] ;
    input \a[1][12] ;
    input \a[1][13] ;
    input \a[1][14] ;
    input \a[1][15] ;
    input \a[2][0] ;
    input \a[2][1] ;
    input \a[2][2] ;
    input \a[2][3] ;
    input \a[2][4] ;
    input \a[2][5] ;
    input \a[2][6] ;
    input \a[2][7] ;
    input \a[2][8] ;
    input \a[2][9] ;
    input \a[2][10] ;
    input \a[2][11] ;
    input \a[2][12] ;
    input \a[2][13] ;
    input \a[2][14] ;
    input \a[2][15] ;
    input \a[3][0] ;
    input \a[3][1] ;
    input \a[3][2] ;
    input \a[3][3] ;
    input \a[3][4] ;
    input \a[3][5] ;
    input \a[3][6] ;
    input \a[3][7] ;
    input \a[3][8] ;
    input \a[3][9] ;
    input \a[3][10] ;
    input \a[3][11] ;
    input \a[3][12] ;
    input \a[3][13] ;
    input \a[3][14] ;
    input \a[3][15] ;
    input \a[4][0] ;
    input \a[4][1] ;
    input \a[4][2] ;
    input \a[4][3] ;
    input \a[4][4] ;
    input \a[4][5] ;
    input \a[4][6] ;
    input \a[4][7] ;
    input \a[4][8] ;
    input \a[4][9] ;
    input \a[4][10] ;
    input \a[4][11] ;
    input \a[4][12] ;
    input \a[4][13] ;
    input \a[4][14] ;
    input \a[4][15] ;
    input \a[5][0] ;
    input \a[5][1] ;
    input \a[5][2] ;
    input \a[5][3] ;
    input \a[5][4] ;
    input \a[5][5] ;
    input \a[5][6] ;
    input \a[5][7] ;
    input \a[5][8] ;
    input \a[5][9] ;
    input \a[5][10] ;
    input \a[5][11] ;
    input \a[5][12] ;
    input \a[5][13] ;
    input \a[5][14] ;
    input \a[5][15] ;
    input \a[6][0] ;
    input \a[6][1] ;
    input \a[6][2] ;
    input \a[6][3] ;
    input \a[6][4] ;
    input \a[6][5] ;
    input \a[6][6] ;
    input \a[6][7] ;
    input \a[6][8] ;
    input \a[6][9] ;
    input \a[6][10] ;
    input \a[6][11] ;
    input \a[6][12] ;
    input \a[6][13] ;
    input \a[6][14] ;
    input \a[6][15] ;
    input \a[7][0] ;
    input \a[7][1] ;
    input \a[7][2] ;
    input \a[7][3] ;
    input \a[7][4] ;
    input \a[7][5] ;
    input \a[7][6] ;
    input \a[7][7] ;
    input \a[7][8] ;
    input \a[7][9] ;
    input \a[7][10] ;
    input \a[7][11] ;
    input \a[7][12] ;
    input \a[7][13] ;
    input \a[7][14] ;
    input \a[7][15] ;
    input \a[8][0] ;
    input \a[8][1] ;
    input \a[8][2] ;
    input \a[8][3] ;
    input \a[8][4] ;
    input \a[8][5] ;
    input \a[8][6] ;
    input \a[8][7] ;
    input \a[8][8] ;
    input \a[8][9] ;
    input \a[8][10] ;
    input \a[8][11] ;
    input \a[8][12] ;
    input \a[8][13] ;
    input \a[8][14] ;
    input \a[8][15] ;
    input \a[9][0] ;
    input \a[9][1] ;
    input \a[9][2] ;
    input \a[9][3] ;
    input \a[9][4] ;
    input \a[9][5] ;
    input \a[9][6] ;
    input \a[9][7] ;
    input \a[9][8] ;
    input \a[9][9] ;
    input \a[9][10] ;
    input \a[9][11] ;
    input \a[9][12] ;
    input \a[9][13] ;
    input \a[9][14] ;
    input \a[9][15] ;
    input \a[10][0] ;
    input \a[10][1] ;
    input \a[10][2] ;
    input \a[10][3] ;
    input \a[10][4] ;
    input \a[10][5] ;
    input \a[10][6] ;
    input \a[10][7] ;
    input \a[10][8] ;
    input \a[10][9] ;
    input \a[10][10] ;
    input \a[10][11] ;
    input \a[10][12] ;
    input \a[10][13] ;
    input \a[10][14] ;
    input \a[10][15] ;
    input \a[11][0] ;
    input \a[11][1] ;
    input \a[11][2] ;
    input \a[11][3] ;
    input \a[11][4] ;
    input \a[11][5] ;
    input \a[11][6] ;
    input \a[11][7] ;
    input \a[11][8] ;
    input \a[11][9] ;
    input \a[11][10] ;
    input \a[11][11] ;
    input \a[11][12] ;
    input \a[11][13] ;
    input \a[11][14] ;
    input \a[11][15] ;
    input \a[12][0] ;
    input \a[12][1] ;
    input \a[12][2] ;
    input \a[12][3] ;
    input \a[12][4] ;
    input \a[12][5] ;
    input \a[12][6] ;
    input \a[12][7] ;
    input \a[12][8] ;
    input \a[12][9] ;
    input \a[12][10] ;
    input \a[12][11] ;
    input \a[12][12] ;
    input \a[12][13] ;
    input \a[12][14] ;
    input \a[12][15] ;
    input \a[13][0] ;
    input \a[13][1] ;
    input \a[13][2] ;
    input \a[13][3] ;
    input \a[13][4] ;
    input \a[13][5] ;
    input \a[13][6] ;
    input \a[13][7] ;
    input \a[13][8] ;
    input \a[13][9] ;
    input \a[13][10] ;
    input \a[13][11] ;
    input \a[13][12] ;
    input \a[13][13] ;
    input \a[13][14] ;
    input \a[13][15] ;
    input \a[14][0] ;
    input \a[14][1] ;
    input \a[14][2] ;
    input \a[14][3] ;
    input \a[14][4] ;
    input \a[14][5] ;
    input \a[14][6] ;
    input \a[14][7] ;
    input \a[14][8] ;
    input \a[14][9] ;
    input \a[14][10] ;
    input \a[14][11] ;
    input \a[14][12] ;
    input \a[14][13] ;
    input \a[14][14] ;
    input \a[14][15] ;
    input \a[15][0] ;
    input \a[15][1] ;
    input \a[15][2] ;
    input \a[15][3] ;
    input \a[15][4] ;
    input \a[15][5] ;
    input \a[15][6] ;
    input \a[15][7] ;
    input \a[15][8] ;
    input \a[15][9] ;
    input \a[15][10] ;
    input \a[15][11] ;
    input \a[15][12] ;
    input \a[15][13] ;
    input \a[15][14] ;
    input \a[15][15] ;
    output \a_sorted[0][0] ;
    reg \a_sorted[0][0] ;
    output \a_sorted[0][1] ;
    reg \a_sorted[0][1] ;
    output \a_sorted[0][2] ;
    reg \a_sorted[0][2] ;
    output \a_sorted[0][3] ;
    reg \a_sorted[0][3] ;
    output \a_sorted[0][4] ;
    reg \a_sorted[0][4] ;
    output \a_sorted[0][5] ;
    reg \a_sorted[0][5] ;
    output \a_sorted[0][6] ;
    reg \a_sorted[0][6] ;
    output \a_sorted[0][7] ;
    reg \a_sorted[0][7] ;
    output \a_sorted[0][8] ;
    reg \a_sorted[0][8] ;
    output \a_sorted[0][9] ;
    reg \a_sorted[0][9] ;
    output \a_sorted[0][10] ;
    reg \a_sorted[0][10] ;
    output \a_sorted[0][11] ;
    reg \a_sorted[0][11] ;
    output \a_sorted[0][12] ;
    reg \a_sorted[0][12] ;
    output \a_sorted[0][13] ;
    reg \a_sorted[0][13] ;
    output \a_sorted[0][14] ;
    reg \a_sorted[0][14] ;
    output \a_sorted[0][15] ;
    reg \a_sorted[0][15] ;
    output \a_sorted[1][0] ;
    reg \a_sorted[1][0] ;
    output \a_sorted[1][1] ;
    reg \a_sorted[1][1] ;
    output \a_sorted[1][2] ;
    reg \a_sorted[1][2] ;
    output \a_sorted[1][3] ;
    reg \a_sorted[1][3] ;
    output \a_sorted[1][4] ;
    reg \a_sorted[1][4] ;
    output \a_sorted[1][5] ;
    reg \a_sorted[1][5] ;
    output \a_sorted[1][6] ;
    reg \a_sorted[1][6] ;
    output \a_sorted[1][7] ;
    reg \a_sorted[1][7] ;
    output \a_sorted[1][8] ;
    reg \a_sorted[1][8] ;
    output \a_sorted[1][9] ;
    reg \a_sorted[1][9] ;
    output \a_sorted[1][10] ;
    reg \a_sorted[1][10] ;
    output \a_sorted[1][11] ;
    reg \a_sorted[1][11] ;
    output \a_sorted[1][12] ;
    reg \a_sorted[1][12] ;
    output \a_sorted[1][13] ;
    reg \a_sorted[1][13] ;
    output \a_sorted[1][14] ;
    reg \a_sorted[1][14] ;
    output \a_sorted[1][15] ;
    reg \a_sorted[1][15] ;
    output \a_sorted[2][0] ;
    reg \a_sorted[2][0] ;
    output \a_sorted[2][1] ;
    reg \a_sorted[2][1] ;
    output \a_sorted[2][2] ;
    reg \a_sorted[2][2] ;
    output \a_sorted[2][3] ;
    reg \a_sorted[2][3] ;
    output \a_sorted[2][4] ;
    reg \a_sorted[2][4] ;
    output \a_sorted[2][5] ;
    reg \a_sorted[2][5] ;
    output \a_sorted[2][6] ;
    reg \a_sorted[2][6] ;
    output \a_sorted[2][7] ;
    reg \a_sorted[2][7] ;
    output \a_sorted[2][8] ;
    reg \a_sorted[2][8] ;
    output \a_sorted[2][9] ;
    reg \a_sorted[2][9] ;
    output \a_sorted[2][10] ;
    reg \a_sorted[2][10] ;
    output \a_sorted[2][11] ;
    reg \a_sorted[2][11] ;
    output \a_sorted[2][12] ;
    reg \a_sorted[2][12] ;
    output \a_sorted[2][13] ;
    reg \a_sorted[2][13] ;
    output \a_sorted[2][14] ;
    reg \a_sorted[2][14] ;
    output \a_sorted[2][15] ;
    reg \a_sorted[2][15] ;
    output \a_sorted[3][0] ;
    reg \a_sorted[3][0] ;
    output \a_sorted[3][1] ;
    reg \a_sorted[3][1] ;
    output \a_sorted[3][2] ;
    reg \a_sorted[3][2] ;
    output \a_sorted[3][3] ;
    reg \a_sorted[3][3] ;
    output \a_sorted[3][4] ;
    reg \a_sorted[3][4] ;
    output \a_sorted[3][5] ;
    reg \a_sorted[3][5] ;
    output \a_sorted[3][6] ;
    reg \a_sorted[3][6] ;
    output \a_sorted[3][7] ;
    reg \a_sorted[3][7] ;
    output \a_sorted[3][8] ;
    reg \a_sorted[3][8] ;
    output \a_sorted[3][9] ;
    reg \a_sorted[3][9] ;
    output \a_sorted[3][10] ;
    reg \a_sorted[3][10] ;
    output \a_sorted[3][11] ;
    reg \a_sorted[3][11] ;
    output \a_sorted[3][12] ;
    reg \a_sorted[3][12] ;
    output \a_sorted[3][13] ;
    reg \a_sorted[3][13] ;
    output \a_sorted[3][14] ;
    reg \a_sorted[3][14] ;
    output \a_sorted[3][15] ;
    reg \a_sorted[3][15] ;
    output \a_sorted[4][0] ;
    reg \a_sorted[4][0] ;
    output \a_sorted[4][1] ;
    reg \a_sorted[4][1] ;
    output \a_sorted[4][2] ;
    reg \a_sorted[4][2] ;
    output \a_sorted[4][3] ;
    reg \a_sorted[4][3] ;
    output \a_sorted[4][4] ;
    reg \a_sorted[4][4] ;
    output \a_sorted[4][5] ;
    reg \a_sorted[4][5] ;
    output \a_sorted[4][6] ;
    reg \a_sorted[4][6] ;
    output \a_sorted[4][7] ;
    reg \a_sorted[4][7] ;
    output \a_sorted[4][8] ;
    reg \a_sorted[4][8] ;
    output \a_sorted[4][9] ;
    reg \a_sorted[4][9] ;
    output \a_sorted[4][10] ;
    reg \a_sorted[4][10] ;
    output \a_sorted[4][11] ;
    reg \a_sorted[4][11] ;
    output \a_sorted[4][12] ;
    reg \a_sorted[4][12] ;
    output \a_sorted[4][13] ;
    reg \a_sorted[4][13] ;
    output \a_sorted[4][14] ;
    reg \a_sorted[4][14] ;
    output \a_sorted[4][15] ;
    reg \a_sorted[4][15] ;
    output \a_sorted[5][0] ;
    reg \a_sorted[5][0] ;
    output \a_sorted[5][1] ;
    reg \a_sorted[5][1] ;
    output \a_sorted[5][2] ;
    reg \a_sorted[5][2] ;
    output \a_sorted[5][3] ;
    reg \a_sorted[5][3] ;
    output \a_sorted[5][4] ;
    reg \a_sorted[5][4] ;
    output \a_sorted[5][5] ;
    reg \a_sorted[5][5] ;
    output \a_sorted[5][6] ;
    reg \a_sorted[5][6] ;
    output \a_sorted[5][7] ;
    reg \a_sorted[5][7] ;
    output \a_sorted[5][8] ;
    reg \a_sorted[5][8] ;
    output \a_sorted[5][9] ;
    reg \a_sorted[5][9] ;
    output \a_sorted[5][10] ;
    reg \a_sorted[5][10] ;
    output \a_sorted[5][11] ;
    reg \a_sorted[5][11] ;
    output \a_sorted[5][12] ;
    reg \a_sorted[5][12] ;
    output \a_sorted[5][13] ;
    reg \a_sorted[5][13] ;
    output \a_sorted[5][14] ;
    reg \a_sorted[5][14] ;
    output \a_sorted[5][15] ;
    reg \a_sorted[5][15] ;
    output \a_sorted[6][0] ;
    reg \a_sorted[6][0] ;
    output \a_sorted[6][1] ;
    reg \a_sorted[6][1] ;
    output \a_sorted[6][2] ;
    reg \a_sorted[6][2] ;
    output \a_sorted[6][3] ;
    reg \a_sorted[6][3] ;
    output \a_sorted[6][4] ;
    reg \a_sorted[6][4] ;
    output \a_sorted[6][5] ;
    reg \a_sorted[6][5] ;
    output \a_sorted[6][6] ;
    reg \a_sorted[6][6] ;
    output \a_sorted[6][7] ;
    reg \a_sorted[6][7] ;
    output \a_sorted[6][8] ;
    reg \a_sorted[6][8] ;
    output \a_sorted[6][9] ;
    reg \a_sorted[6][9] ;
    output \a_sorted[6][10] ;
    reg \a_sorted[6][10] ;
    output \a_sorted[6][11] ;
    reg \a_sorted[6][11] ;
    output \a_sorted[6][12] ;
    reg \a_sorted[6][12] ;
    output \a_sorted[6][13] ;
    reg \a_sorted[6][13] ;
    output \a_sorted[6][14] ;
    reg \a_sorted[6][14] ;
    output \a_sorted[6][15] ;
    reg \a_sorted[6][15] ;
    output \a_sorted[7][0] ;
    reg \a_sorted[7][0] ;
    output \a_sorted[7][1] ;
    reg \a_sorted[7][1] ;
    output \a_sorted[7][2] ;
    reg \a_sorted[7][2] ;
    output \a_sorted[7][3] ;
    reg \a_sorted[7][3] ;
    output \a_sorted[7][4] ;
    reg \a_sorted[7][4] ;
    output \a_sorted[7][5] ;
    reg \a_sorted[7][5] ;
    output \a_sorted[7][6] ;
    reg \a_sorted[7][6] ;
    output \a_sorted[7][7] ;
    reg \a_sorted[7][7] ;
    output \a_sorted[7][8] ;
    reg \a_sorted[7][8] ;
    output \a_sorted[7][9] ;
    reg \a_sorted[7][9] ;
    output \a_sorted[7][10] ;
    reg \a_sorted[7][10] ;
    output \a_sorted[7][11] ;
    reg \a_sorted[7][11] ;
    output \a_sorted[7][12] ;
    reg \a_sorted[7][12] ;
    output \a_sorted[7][13] ;
    reg \a_sorted[7][13] ;
    output \a_sorted[7][14] ;
    reg \a_sorted[7][14] ;
    output \a_sorted[7][15] ;
    reg \a_sorted[7][15] ;
    output \a_sorted[8][0] ;
    reg \a_sorted[8][0] ;
    output \a_sorted[8][1] ;
    reg \a_sorted[8][1] ;
    output \a_sorted[8][2] ;
    reg \a_sorted[8][2] ;
    output \a_sorted[8][3] ;
    reg \a_sorted[8][3] ;
    output \a_sorted[8][4] ;
    reg \a_sorted[8][4] ;
    output \a_sorted[8][5] ;
    reg \a_sorted[8][5] ;
    output \a_sorted[8][6] ;
    reg \a_sorted[8][6] ;
    output \a_sorted[8][7] ;
    reg \a_sorted[8][7] ;
    output \a_sorted[8][8] ;
    reg \a_sorted[8][8] ;
    output \a_sorted[8][9] ;
    reg \a_sorted[8][9] ;
    output \a_sorted[8][10] ;
    reg \a_sorted[8][10] ;
    output \a_sorted[8][11] ;
    reg \a_sorted[8][11] ;
    output \a_sorted[8][12] ;
    reg \a_sorted[8][12] ;
    output \a_sorted[8][13] ;
    reg \a_sorted[8][13] ;
    output \a_sorted[8][14] ;
    reg \a_sorted[8][14] ;
    output \a_sorted[8][15] ;
    reg \a_sorted[8][15] ;
    output \a_sorted[9][0] ;
    reg \a_sorted[9][0] ;
    output \a_sorted[9][1] ;
    reg \a_sorted[9][1] ;
    output \a_sorted[9][2] ;
    reg \a_sorted[9][2] ;
    output \a_sorted[9][3] ;
    reg \a_sorted[9][3] ;
    output \a_sorted[9][4] ;
    reg \a_sorted[9][4] ;
    output \a_sorted[9][5] ;
    reg \a_sorted[9][5] ;
    output \a_sorted[9][6] ;
    reg \a_sorted[9][6] ;
    output \a_sorted[9][7] ;
    reg \a_sorted[9][7] ;
    output \a_sorted[9][8] ;
    reg \a_sorted[9][8] ;
    output \a_sorted[9][9] ;
    reg \a_sorted[9][9] ;
    output \a_sorted[9][10] ;
    reg \a_sorted[9][10] ;
    output \a_sorted[9][11] ;
    reg \a_sorted[9][11] ;
    output \a_sorted[9][12] ;
    reg \a_sorted[9][12] ;
    output \a_sorted[9][13] ;
    reg \a_sorted[9][13] ;
    output \a_sorted[9][14] ;
    reg \a_sorted[9][14] ;
    output \a_sorted[9][15] ;
    reg \a_sorted[9][15] ;
    output \a_sorted[10][0] ;
    reg \a_sorted[10][0] ;
    output \a_sorted[10][1] ;
    reg \a_sorted[10][1] ;
    output \a_sorted[10][2] ;
    reg \a_sorted[10][2] ;
    output \a_sorted[10][3] ;
    reg \a_sorted[10][3] ;
    output \a_sorted[10][4] ;
    reg \a_sorted[10][4] ;
    output \a_sorted[10][5] ;
    reg \a_sorted[10][5] ;
    output \a_sorted[10][6] ;
    reg \a_sorted[10][6] ;
    output \a_sorted[10][7] ;
    reg \a_sorted[10][7] ;
    output \a_sorted[10][8] ;
    reg \a_sorted[10][8] ;
    output \a_sorted[10][9] ;
    reg \a_sorted[10][9] ;
    output \a_sorted[10][10] ;
    reg \a_sorted[10][10] ;
    output \a_sorted[10][11] ;
    reg \a_sorted[10][11] ;
    output \a_sorted[10][12] ;
    reg \a_sorted[10][12] ;
    output \a_sorted[10][13] ;
    reg \a_sorted[10][13] ;
    output \a_sorted[10][14] ;
    reg \a_sorted[10][14] ;
    output \a_sorted[10][15] ;
    reg \a_sorted[10][15] ;
    output \a_sorted[11][0] ;
    reg \a_sorted[11][0] ;
    output \a_sorted[11][1] ;
    reg \a_sorted[11][1] ;
    output \a_sorted[11][2] ;
    reg \a_sorted[11][2] ;
    output \a_sorted[11][3] ;
    reg \a_sorted[11][3] ;
    output \a_sorted[11][4] ;
    reg \a_sorted[11][4] ;
    output \a_sorted[11][5] ;
    reg \a_sorted[11][5] ;
    output \a_sorted[11][6] ;
    reg \a_sorted[11][6] ;
    output \a_sorted[11][7] ;
    reg \a_sorted[11][7] ;
    output \a_sorted[11][8] ;
    reg \a_sorted[11][8] ;
    output \a_sorted[11][9] ;
    reg \a_sorted[11][9] ;
    output \a_sorted[11][10] ;
    reg \a_sorted[11][10] ;
    output \a_sorted[11][11] ;
    reg \a_sorted[11][11] ;
    output \a_sorted[11][12] ;
    reg \a_sorted[11][12] ;
    output \a_sorted[11][13] ;
    reg \a_sorted[11][13] ;
    output \a_sorted[11][14] ;
    reg \a_sorted[11][14] ;
    output \a_sorted[11][15] ;
    reg \a_sorted[11][15] ;
    output \a_sorted[12][0] ;
    reg \a_sorted[12][0] ;
    output \a_sorted[12][1] ;
    reg \a_sorted[12][1] ;
    output \a_sorted[12][2] ;
    reg \a_sorted[12][2] ;
    output \a_sorted[12][3] ;
    reg \a_sorted[12][3] ;
    output \a_sorted[12][4] ;
    reg \a_sorted[12][4] ;
    output \a_sorted[12][5] ;
    reg \a_sorted[12][5] ;
    output \a_sorted[12][6] ;
    reg \a_sorted[12][6] ;
    output \a_sorted[12][7] ;
    reg \a_sorted[12][7] ;
    output \a_sorted[12][8] ;
    reg \a_sorted[12][8] ;
    output \a_sorted[12][9] ;
    reg \a_sorted[12][9] ;
    output \a_sorted[12][10] ;
    reg \a_sorted[12][10] ;
    output \a_sorted[12][11] ;
    reg \a_sorted[12][11] ;
    output \a_sorted[12][12] ;
    reg \a_sorted[12][12] ;
    output \a_sorted[12][13] ;
    reg \a_sorted[12][13] ;
    output \a_sorted[12][14] ;
    reg \a_sorted[12][14] ;
    output \a_sorted[12][15] ;
    reg \a_sorted[12][15] ;
    output \a_sorted[13][0] ;
    reg \a_sorted[13][0] ;
    output \a_sorted[13][1] ;
    reg \a_sorted[13][1] ;
    output \a_sorted[13][2] ;
    reg \a_sorted[13][2] ;
    output \a_sorted[13][3] ;
    reg \a_sorted[13][3] ;
    output \a_sorted[13][4] ;
    reg \a_sorted[13][4] ;
    output \a_sorted[13][5] ;
    reg \a_sorted[13][5] ;
    output \a_sorted[13][6] ;
    reg \a_sorted[13][6] ;
    output \a_sorted[13][7] ;
    reg \a_sorted[13][7] ;
    output \a_sorted[13][8] ;
    reg \a_sorted[13][8] ;
    output \a_sorted[13][9] ;
    reg \a_sorted[13][9] ;
    output \a_sorted[13][10] ;
    reg \a_sorted[13][10] ;
    output \a_sorted[13][11] ;
    reg \a_sorted[13][11] ;
    output \a_sorted[13][12] ;
    reg \a_sorted[13][12] ;
    output \a_sorted[13][13] ;
    reg \a_sorted[13][13] ;
    output \a_sorted[13][14] ;
    reg \a_sorted[13][14] ;
    output \a_sorted[13][15] ;
    reg \a_sorted[13][15] ;
    output \a_sorted[14][0] ;
    reg \a_sorted[14][0] ;
    output \a_sorted[14][1] ;
    reg \a_sorted[14][1] ;
    output \a_sorted[14][2] ;
    reg \a_sorted[14][2] ;
    output \a_sorted[14][3] ;
    reg \a_sorted[14][3] ;
    output \a_sorted[14][4] ;
    reg \a_sorted[14][4] ;
    output \a_sorted[14][5] ;
    reg \a_sorted[14][5] ;
    output \a_sorted[14][6] ;
    reg \a_sorted[14][6] ;
    output \a_sorted[14][7] ;
    reg \a_sorted[14][7] ;
    output \a_sorted[14][8] ;
    reg \a_sorted[14][8] ;
    output \a_sorted[14][9] ;
    reg \a_sorted[14][9] ;
    output \a_sorted[14][10] ;
    reg \a_sorted[14][10] ;
    output \a_sorted[14][11] ;
    reg \a_sorted[14][11] ;
    output \a_sorted[14][12] ;
    reg \a_sorted[14][12] ;
    output \a_sorted[14][13] ;
    reg \a_sorted[14][13] ;
    output \a_sorted[14][14] ;
    reg \a_sorted[14][14] ;
    output \a_sorted[14][15] ;
    reg \a_sorted[14][15] ;
    output \a_sorted[15][0] ;
    reg \a_sorted[15][0] ;
    output \a_sorted[15][1] ;
    reg \a_sorted[15][1] ;
    output \a_sorted[15][2] ;
    reg \a_sorted[15][2] ;
    output \a_sorted[15][3] ;
    reg \a_sorted[15][3] ;
    output \a_sorted[15][4] ;
    reg \a_sorted[15][4] ;
    output \a_sorted[15][5] ;
    reg \a_sorted[15][5] ;
    output \a_sorted[15][6] ;
    reg \a_sorted[15][6] ;
    output \a_sorted[15][7] ;
    reg \a_sorted[15][7] ;
    output \a_sorted[15][8] ;
    reg \a_sorted[15][8] ;
    output \a_sorted[15][9] ;
    reg \a_sorted[15][9] ;
    output \a_sorted[15][10] ;
    reg \a_sorted[15][10] ;
    output \a_sorted[15][11] ;
    reg \a_sorted[15][11] ;
    output \a_sorted[15][12] ;
    reg \a_sorted[15][12] ;
    output \a_sorted[15][13] ;
    reg \a_sorted[15][13] ;
    output \a_sorted[15][14] ;
    reg \a_sorted[15][14] ;
    output \a_sorted[15][15] ;
    reg \a_sorted[15][15] ;
    wire \a_sorted[0][0]_ns ;
    wire \a_sorted[0][1]_ns ;
    wire \a_sorted[0][2]_ns ;
    wire \a_sorted[0][3]_ns ;
    wire \a_sorted[0][4]_ns ;
    wire \a_sorted[0][5]_ns ;
    wire \a_sorted[0][6]_ns ;
    wire \a_sorted[0][7]_ns ;
    wire \a_sorted[0][8]_ns ;
    wire \a_sorted[0][9]_ns ;
    wire \a_sorted[0][10]_ns ;
    wire \a_sorted[0][11]_ns ;
    wire \a_sorted[0][12]_ns ;
    wire \a_sorted[0][13]_ns ;
    wire \a_sorted[0][14]_ns ;
    wire \a_sorted[0][15]_ns ;
    wire \a_sorted[1][0]_ns ;
    wire \a_sorted[1][1]_ns ;
    wire \a_sorted[1][2]_ns ;
    wire \a_sorted[1][3]_ns ;
    wire \a_sorted[1][4]_ns ;
    wire \a_sorted[1][5]_ns ;
    wire \a_sorted[1][6]_ns ;
    wire \a_sorted[1][7]_ns ;
    wire \a_sorted[1][8]_ns ;
    wire \a_sorted[1][9]_ns ;
    wire \a_sorted[1][10]_ns ;
    wire \a_sorted[1][11]_ns ;
    wire \a_sorted[1][12]_ns ;
    wire \a_sorted[1][13]_ns ;
    wire \a_sorted[1][14]_ns ;
    wire \a_sorted[1][15]_ns ;
    wire \a_sorted[2][0]_ns ;
    wire \a_sorted[2][1]_ns ;
    wire \a_sorted[2][2]_ns ;
    wire \a_sorted[2][3]_ns ;
    wire \a_sorted[2][4]_ns ;
    wire \a_sorted[2][5]_ns ;
    wire \a_sorted[2][6]_ns ;
    wire \a_sorted[2][7]_ns ;
    wire \a_sorted[2][8]_ns ;
    wire \a_sorted[2][9]_ns ;
    wire \a_sorted[2][10]_ns ;
    wire \a_sorted[2][11]_ns ;
    wire \a_sorted[2][12]_ns ;
    wire \a_sorted[2][13]_ns ;
    wire \a_sorted[2][14]_ns ;
    wire \a_sorted[2][15]_ns ;
    wire \a_sorted[3][0]_ns ;
    wire \a_sorted[3][1]_ns ;
    wire \a_sorted[3][2]_ns ;
    wire \a_sorted[3][3]_ns ;
    wire \a_sorted[3][4]_ns ;
    wire \a_sorted[3][5]_ns ;
    wire \a_sorted[3][6]_ns ;
    wire \a_sorted[3][7]_ns ;
    wire \a_sorted[3][8]_ns ;
    wire \a_sorted[3][9]_ns ;
    wire \a_sorted[3][10]_ns ;
    wire \a_sorted[3][11]_ns ;
    wire \a_sorted[3][12]_ns ;
    wire \a_sorted[3][13]_ns ;
    wire \a_sorted[3][14]_ns ;
    wire \a_sorted[3][15]_ns ;
    wire \a_sorted[4][0]_ns ;
    wire \a_sorted[4][1]_ns ;
    wire \a_sorted[4][2]_ns ;
    wire \a_sorted[4][3]_ns ;
    wire \a_sorted[4][4]_ns ;
    wire \a_sorted[4][5]_ns ;
    wire \a_sorted[4][6]_ns ;
    wire \a_sorted[4][7]_ns ;
    wire \a_sorted[4][8]_ns ;
    wire \a_sorted[4][9]_ns ;
    wire \a_sorted[4][10]_ns ;
    wire \a_sorted[4][11]_ns ;
    wire \a_sorted[4][12]_ns ;
    wire \a_sorted[4][13]_ns ;
    wire \a_sorted[4][14]_ns ;
    wire \a_sorted[4][15]_ns ;
    wire \a_sorted[5][0]_ns ;
    wire \a_sorted[5][1]_ns ;
    wire \a_sorted[5][2]_ns ;
    wire \a_sorted[5][3]_ns ;
    wire \a_sorted[5][4]_ns ;
    wire \a_sorted[5][5]_ns ;
    wire \a_sorted[5][6]_ns ;
    wire \a_sorted[5][7]_ns ;
    wire \a_sorted[5][8]_ns ;
    wire \a_sorted[5][9]_ns ;
    wire \a_sorted[5][10]_ns ;
    wire \a_sorted[5][11]_ns ;
    wire \a_sorted[5][12]_ns ;
    wire \a_sorted[5][13]_ns ;
    wire \a_sorted[5][14]_ns ;
    wire \a_sorted[5][15]_ns ;
    wire \a_sorted[6][0]_ns ;
    wire \a_sorted[6][1]_ns ;
    wire \a_sorted[6][2]_ns ;
    wire \a_sorted[6][3]_ns ;
    wire \a_sorted[6][4]_ns ;
    wire \a_sorted[6][5]_ns ;
    wire \a_sorted[6][6]_ns ;
    wire \a_sorted[6][7]_ns ;
    wire \a_sorted[6][8]_ns ;
    wire \a_sorted[6][9]_ns ;
    wire \a_sorted[6][10]_ns ;
    wire \a_sorted[6][11]_ns ;
    wire \a_sorted[6][12]_ns ;
    wire \a_sorted[6][13]_ns ;
    wire \a_sorted[6][14]_ns ;
    wire \a_sorted[6][15]_ns ;
    wire \a_sorted[7][0]_ns ;
    wire \a_sorted[7][1]_ns ;
    wire \a_sorted[7][2]_ns ;
    wire \a_sorted[7][3]_ns ;
    wire \a_sorted[7][4]_ns ;
    wire \a_sorted[7][5]_ns ;
    wire \a_sorted[7][6]_ns ;
    wire \a_sorted[7][7]_ns ;
    wire \a_sorted[7][8]_ns ;
    wire \a_sorted[7][9]_ns ;
    wire \a_sorted[7][10]_ns ;
    wire \a_sorted[7][11]_ns ;
    wire \a_sorted[7][12]_ns ;
    wire \a_sorted[7][13]_ns ;
    wire \a_sorted[7][14]_ns ;
    wire \a_sorted[7][15]_ns ;
    wire \a_sorted[8][0]_ns ;
    wire \a_sorted[8][1]_ns ;
    wire \a_sorted[8][2]_ns ;
    wire \a_sorted[8][3]_ns ;
    wire \a_sorted[8][4]_ns ;
    wire \a_sorted[8][5]_ns ;
    wire \a_sorted[8][6]_ns ;
    wire \a_sorted[8][7]_ns ;
    wire \a_sorted[8][8]_ns ;
    wire \a_sorted[8][9]_ns ;
    wire \a_sorted[8][10]_ns ;
    wire \a_sorted[8][11]_ns ;
    wire \a_sorted[8][12]_ns ;
    wire \a_sorted[8][13]_ns ;
    wire \a_sorted[8][14]_ns ;
    wire \a_sorted[8][15]_ns ;
    wire \a_sorted[9][0]_ns ;
    wire \a_sorted[9][1]_ns ;
    wire \a_sorted[9][2]_ns ;
    wire \a_sorted[9][3]_ns ;
    wire \a_sorted[9][4]_ns ;
    wire \a_sorted[9][5]_ns ;
    wire \a_sorted[9][6]_ns ;
    wire \a_sorted[9][7]_ns ;
    wire \a_sorted[9][8]_ns ;
    wire \a_sorted[9][9]_ns ;
    wire \a_sorted[9][10]_ns ;
    wire \a_sorted[9][11]_ns ;
    wire \a_sorted[9][12]_ns ;
    wire \a_sorted[9][13]_ns ;
    wire \a_sorted[9][14]_ns ;
    wire \a_sorted[9][15]_ns ;
    wire \a_sorted[10][0]_ns ;
    wire \a_sorted[10][1]_ns ;
    wire \a_sorted[10][2]_ns ;
    wire \a_sorted[10][3]_ns ;
    wire \a_sorted[10][4]_ns ;
    wire \a_sorted[10][5]_ns ;
    wire \a_sorted[10][6]_ns ;
    wire \a_sorted[10][7]_ns ;
    wire \a_sorted[10][8]_ns ;
    wire \a_sorted[10][9]_ns ;
    wire \a_sorted[10][10]_ns ;
    wire \a_sorted[10][11]_ns ;
    wire \a_sorted[10][12]_ns ;
    wire \a_sorted[10][13]_ns ;
    wire \a_sorted[10][14]_ns ;
    wire \a_sorted[10][15]_ns ;
    wire \a_sorted[11][0]_ns ;
    wire \a_sorted[11][1]_ns ;
    wire \a_sorted[11][2]_ns ;
    wire \a_sorted[11][3]_ns ;
    wire \a_sorted[11][4]_ns ;
    wire \a_sorted[11][5]_ns ;
    wire \a_sorted[11][6]_ns ;
    wire \a_sorted[11][7]_ns ;
    wire \a_sorted[11][8]_ns ;
    wire \a_sorted[11][9]_ns ;
    wire \a_sorted[11][10]_ns ;
    wire \a_sorted[11][11]_ns ;
    wire \a_sorted[11][12]_ns ;
    wire \a_sorted[11][13]_ns ;
    wire \a_sorted[11][14]_ns ;
    wire \a_sorted[11][15]_ns ;
    wire \a_sorted[12][0]_ns ;
    wire \a_sorted[12][1]_ns ;
    wire \a_sorted[12][2]_ns ;
    wire \a_sorted[12][3]_ns ;
    wire \a_sorted[12][4]_ns ;
    wire \a_sorted[12][5]_ns ;
    wire \a_sorted[12][6]_ns ;
    wire \a_sorted[12][7]_ns ;
    wire \a_sorted[12][8]_ns ;
    wire \a_sorted[12][9]_ns ;
    wire \a_sorted[12][10]_ns ;
    wire \a_sorted[12][11]_ns ;
    wire \a_sorted[12][12]_ns ;
    wire \a_sorted[12][13]_ns ;
    wire \a_sorted[12][14]_ns ;
    wire \a_sorted[12][15]_ns ;
    wire \a_sorted[13][0]_ns ;
    wire \a_sorted[13][1]_ns ;
    wire \a_sorted[13][2]_ns ;
    wire \a_sorted[13][3]_ns ;
    wire \a_sorted[13][4]_ns ;
    wire \a_sorted[13][5]_ns ;
    wire \a_sorted[13][6]_ns ;
    wire \a_sorted[13][7]_ns ;
    wire \a_sorted[13][8]_ns ;
    wire \a_sorted[13][9]_ns ;
    wire \a_sorted[13][10]_ns ;
    wire \a_sorted[13][11]_ns ;
    wire \a_sorted[13][12]_ns ;
    wire \a_sorted[13][13]_ns ;
    wire \a_sorted[13][14]_ns ;
    wire \a_sorted[13][15]_ns ;
    wire \a_sorted[14][0]_ns ;
    wire \a_sorted[14][1]_ns ;
    wire \a_sorted[14][2]_ns ;
    wire \a_sorted[14][3]_ns ;
    wire \a_sorted[14][4]_ns ;
    wire \a_sorted[14][5]_ns ;
    wire \a_sorted[14][6]_ns ;
    wire \a_sorted[14][7]_ns ;
    wire \a_sorted[14][8]_ns ;
    wire \a_sorted[14][9]_ns ;
    wire \a_sorted[14][10]_ns ;
    wire \a_sorted[14][11]_ns ;
    wire \a_sorted[14][12]_ns ;
    wire \a_sorted[14][13]_ns ;
    wire \a_sorted[14][14]_ns ;
    wire \a_sorted[14][15]_ns ;
    wire \a_sorted[15][0]_ns ;
    wire \a_sorted[15][1]_ns ;
    wire \a_sorted[15][2]_ns ;
    wire \a_sorted[15][3]_ns ;
    wire \a_sorted[15][4]_ns ;
    wire \a_sorted[15][5]_ns ;
    wire \a_sorted[15][6]_ns ;
    wire \a_sorted[15][7]_ns ;
    wire \a_sorted[15][8]_ns ;
    wire \a_sorted[15][9]_ns ;
    wire \a_sorted[15][10]_ns ;
    wire \a_sorted[15][11]_ns ;
    wire \a_sorted[15][12]_ns ;
    wire \a_sorted[15][13]_ns ;
    wire \a_sorted[15][14]_ns ;
    wire \a_sorted[15][15]_ns ;
    wire _0;
    wire _1;
    wire _2;
    wire _3;
    wire _4;
    wire _5;
    wire _6;
    wire _7;
    wire _8;
    wire _9;
    wire _10;
    wire _11;
    wire _12;
    wire _13;
    wire _14;
    wire _15;
    wire _16;
    wire _17;
    wire _18;
    wire _19;
    wire _20;
    wire _21;
    wire _22;
    wire _23;
    wire _24;
    wire _25;
    wire _26;
    wire _27;
    wire _28;
    wire _29;
    wire _30;
    wire _31;
    wire _32;
    wire _33;
    wire _34;
    wire _35;
    wire _36;
    wire _37;
    wire _38;
    wire _39;
    wire _40;
    wire _41;
    wire _42;
    wire _43;
    wire _44;
    wire _45;
    wire _46;
    wire _47;
    wire _48;
    wire _49;
    wire _50;
    wire _51;
    wire _52;
    wire _53;
    wire _54;
    wire _55;
    wire _56;
    wire _57;
    wire _58;
    wire _59;
    wire _60;
    wire _61;
    wire _62;
    wire _63;
    wire _64;
    wire _65;
    wire _66;
    wire _67;
    wire _68;
    wire _69;
    wire _70;
    wire _71;
    wire _72;
    wire _73;
    wire _74;
    wire _75;
    wire _76;
    wire _77;
    wire _78;
    wire _79;
    wire _80;
    wire _81;
    wire _82;
    wire _83;
    wire _84;
    wire _85;
    wire _86;
    wire _87;
    wire _88;
    wire _89;
    wire _90;
    wire _91;
    wire _92;
    wire _93;
    wire _94;
    wire _95;
    wire _96;
    wire _97;
    wire _98;
    wire _99;
    wire _100;
    wire _101;
    wire _102;
    wire _103;
    wire _104;
    wire _105;
    wire _106;
    wire _107;
    wire _108;
    wire _109;
    wire _110;
    wire _111;
    wire _112;
    wire _113;
    wire _114;
    wire _115;
    wire _116;
    wire _117;
    wire _118;
    wire _119;
    wire _120;
    wire _121;
    wire _122;
    wire _123;
    wire _124;
    wire _125;
    wire _126;
    wire _127;
    wire _128;
    wire _129;
    wire _130;
    wire _131;
    wire _132;
    wire _133;
    wire _134;
    wire _135;
    wire _136;
    wire _137;
    wire _138;
    wire _139;
    wire _140;
    wire _141;
    wire _142;
    wire _143;
    wire _144;
    wire _145;
    wire _146;
    wire _147;
    wire _148;
    wire _149;
    wire _150;
    wire _151;
    wire _152;
    wire _153;
    wire _154;
    wire _155;
    wire _156;
    wire _157;
    wire _158;
    wire _159;
    wire _160;
    wire _161;
    wire _162;
    wire _163;
    wire _164;
    wire _165;
    wire _166;
    wire _167;
    wire _168;
    wire _169;
    wire _170;
    wire _171;
    wire _172;
    wire _173;
    wire _174;
    wire _175;
    wire _176;
    wire _177;
    wire _178;
    wire _179;
    wire _180;
    wire _181;
    wire _182;
    wire _183;
    wire _184;
    wire _185;
    wire _186;
    wire _187;
    wire _188;
    wire _189;
    wire _190;
    wire _191;
    wire _192;
    wire _193;
    wire _194;
    wire _195;
    wire _196;
    wire _197;
    wire _198;
    wire _199;
    wire _200;
    wire _201;
    wire _202;
    wire _203;
    wire _204;
    wire _205;
    wire _206;
    wire _207;
    wire _208;
    wire _209;
    wire _210;
    wire _211;
    wire _212;
    wire _213;
    wire _214;
    wire _215;
    wire _216;
    wire _217;
    wire _218;
    wire _219;
    wire _220;
    wire _221;
    wire _222;
    wire _223;
    wire _224;
    wire _225;
    wire _226;
    wire _227;
    wire _228;
    wire _229;
    wire _230;
    wire _231;
    wire _232;
    wire _233;
    wire _234;
    wire _235;
    wire _236;
    wire _237;
    wire _238;
    wire _239;
    wire _240;
    wire _241;
    wire _242;
    wire _243;
    wire _244;
    wire _245;
    wire _246;
    wire _247;
    wire _248;
    wire _249;
    wire _250;
    wire _251;
    wire _252;
    wire _253;
    wire _254;
    wire _255;
    wire _289;
    wire _290;
    wire _291;
    wire _292;
    wire _293;
    wire _294;
    wire _295;
    wire _296;
    wire _297;
    wire _298;
    wire _299;
    wire _300;
    wire _301;
    wire _302;
    wire _303;
    wire _304;
    wire _305;
    wire _306;
    wire _307;
    wire _308;
    wire _309;
    wire _310;
    wire _311;
    wire _312;
    wire _313;
    wire _314;
    wire _315;
    wire _316;
    wire _317;
    wire _318;
    wire _319;
    wire _320;
    wire _354;
    wire _355;
    wire _356;
    wire _357;
    wire _358;
    wire _359;
    wire _360;
    wire _361;
    wire _362;
    wire _363;
    wire _364;
    wire _365;
    wire _366;
    wire _367;
    wire _368;
    wire _369;
    wire _370;
    wire _371;
    wire _372;
    wire _373;
    wire _374;
    wire _375;
    wire _376;
    wire _377;
    wire _378;
    wire _379;
    wire _380;
    wire _381;
    wire _382;
    wire _383;
    wire _384;
    wire _385;
    wire _419;
    wire _420;
    wire _421;
    wire _422;
    wire _423;
    wire _424;
    wire _425;
    wire _426;
    wire _427;
    wire _428;
    wire _429;
    wire _430;
    wire _431;
    wire _432;
    wire _433;
    wire _434;
    wire _435;
    wire _436;
    wire _437;
    wire _438;
    wire _439;
    wire _440;
    wire _441;
    wire _442;
    wire _443;
    wire _444;
    wire _445;
    wire _446;
    wire _447;
    wire _448;
    wire _449;
    wire _450;
    wire _484;
    wire _485;
    wire _486;
    wire _487;
    wire _488;
    wire _489;
    wire _490;
    wire _491;
    wire _492;
    wire _493;
    wire _494;
    wire _495;
    wire _496;
    wire _497;
    wire _498;
    wire _499;
    wire _500;
    wire _501;
    wire _502;
    wire _503;
    wire _504;
    wire _505;
    wire _506;
    wire _507;
    wire _508;
    wire _509;
    wire _510;
    wire _511;
    wire _512;
    wire _513;
    wire _514;
    wire _515;
    wire _549;
    wire _550;
    wire _551;
    wire _552;
    wire _553;
    wire _554;
    wire _555;
    wire _556;
    wire _557;
    wire _558;
    wire _559;
    wire _560;
    wire _561;
    wire _562;
    wire _563;
    wire _564;
    wire _565;
    wire _566;
    wire _567;
    wire _568;
    wire _569;
    wire _570;
    wire _571;
    wire _572;
    wire _573;
    wire _574;
    wire _575;
    wire _576;
    wire _577;
    wire _578;
    wire _579;
    wire _580;
    wire _614;
    wire _615;
    wire _616;
    wire _617;
    wire _618;
    wire _619;
    wire _620;
    wire _621;
    wire _622;
    wire _623;
    wire _624;
    wire _625;
    wire _626;
    wire _627;
    wire _628;
    wire _629;
    wire _630;
    wire _631;
    wire _632;
    wire _633;
    wire _634;
    wire _635;
    wire _636;
    wire _637;
    wire _638;
    wire _639;
    wire _640;
    wire _641;
    wire _642;
    wire _643;
    wire _644;
    wire _645;
    wire _679;
    wire _680;
    wire _681;
    wire _682;
    wire _683;
    wire _684;
    wire _685;
    wire _686;
    wire _687;
    wire _688;
    wire _689;
    wire _690;
    wire _691;
    wire _692;
    wire _693;
    wire _694;
    wire _695;
    wire _696;
    wire _697;
    wire _698;
    wire _699;
    wire _700;
    wire _701;
    wire _702;
    wire _703;
    wire _704;
    wire _705;
    wire _706;
    wire _707;
    wire _708;
    wire _709;
    wire _710;
    wire _744;
    wire _745;
    wire _746;
    wire _747;
    wire _748;
    wire _749;
    wire _750;
    wire _751;
    wire _752;
    wire _753;
    wire _754;
    wire _755;
    wire _756;
    wire _757;
    wire _758;
    wire _759;
    wire _760;
    wire _761;
    wire _762;
    wire _763;
    wire _764;
    wire _765;
    wire _766;
    wire _767;
    wire _768;
    wire _769;
    wire _770;
    wire _771;
    wire _772;
    wire _773;
    wire _774;
    wire _775;
    wire _809;
    wire _810;
    wire _811;
    wire _812;
    wire _813;
    wire _814;
    wire _815;
    wire _816;
    wire _817;
    wire _818;
    wire _819;
    wire _820;
    wire _821;
    wire _822;
    wire _823;
    wire _824;
    wire _825;
    wire _826;
    wire _827;
    wire _828;
    wire _829;
    wire _830;
    wire _831;
    wire _832;
    wire _833;
    wire _834;
    wire _835;
    wire _836;
    wire _837;
    wire _838;
    wire _839;
    wire _840;
    wire _874;
    wire _875;
    wire _876;
    wire _877;
    wire _878;
    wire _879;
    wire _880;
    wire _881;
    wire _882;
    wire _883;
    wire _884;
    wire _885;
    wire _886;
    wire _887;
    wire _888;
    wire _889;
    wire _890;
    wire _891;
    wire _892;
    wire _893;
    wire _894;
    wire _895;
    wire _896;
    wire _897;
    wire _898;
    wire _899;
    wire _900;
    wire _901;
    wire _902;
    wire _903;
    wire _904;
    wire _905;
    wire _939;
    wire _940;
    wire _941;
    wire _942;
    wire _943;
    wire _944;
    wire _945;
    wire _946;
    wire _947;
    wire _948;
    wire _949;
    wire _950;
    wire _951;
    wire _952;
    wire _953;
    wire _954;
    wire _955;
    wire _956;
    wire _957;
    wire _958;
    wire _959;
    wire _960;
    wire _961;
    wire _962;
    wire _963;
    wire _964;
    wire _965;
    wire _966;
    wire _967;
    wire _968;
    wire _969;
    wire _970;
    wire _1004;
    wire _1005;
    wire _1006;
    wire _1007;
    wire _1008;
    wire _1009;
    wire _1010;
    wire _1011;
    wire _1012;
    wire _1013;
    wire _1014;
    wire _1015;
    wire _1016;
    wire _1017;
    wire _1018;
    wire _1019;
    wire _1020;
    wire _1021;
    wire _1022;
    wire _1023;
    wire _1024;
    wire _1025;
    wire _1026;
    wire _1027;
    wire _1028;
    wire _1029;
    wire _1030;
    wire _1031;
    wire _1032;
    wire _1033;
    wire _1034;
    wire _1035;
    wire _1069;
    wire _1070;
    wire _1071;
    wire _1072;
    wire _1073;
    wire _1074;
    wire _1075;
    wire _1076;
    wire _1077;
    wire _1078;
    wire _1079;
    wire _1080;
    wire _1081;
    wire _1082;
    wire _1083;
    wire _1084;
    wire _1085;
    wire _1086;
    wire _1087;
    wire _1088;
    wire _1089;
    wire _1090;
    wire _1091;
    wire _1092;
    wire _1093;
    wire _1094;
    wire _1095;
    wire _1096;
    wire _1097;
    wire _1098;
    wire _1099;
    wire _1100;
    wire _1134;
    wire _1135;
    wire _1136;
    wire _1137;
    wire _1138;
    wire _1139;
    wire _1140;
    wire _1141;
    wire _1142;
    wire _1143;
    wire _1144;
    wire _1145;
    wire _1146;
    wire _1147;
    wire _1148;
    wire _1149;
    wire _1150;
    wire _1151;
    wire _1152;
    wire _1153;
    wire _1154;
    wire _1155;
    wire _1156;
    wire _1157;
    wire _1158;
    wire _1159;
    wire _1160;
    wire _1161;
    wire _1162;
    wire _1163;
    wire _1164;
    wire _1165;
    wire _1199;
    wire _1200;
    wire _1201;
    wire _1202;
    wire _1203;
    wire _1204;
    wire _1205;
    wire _1206;
    wire _1207;
    wire _1208;
    wire _1209;
    wire _1210;
    wire _1211;
    wire _1212;
    wire _1213;
    wire _1214;
    wire _1215;
    wire _1216;
    wire _1217;
    wire _1218;
    wire _1219;
    wire _1220;
    wire _1221;
    wire _1222;
    wire _1223;
    wire _1224;
    wire _1225;
    wire _1226;
    wire _1227;
    wire _1228;
    wire _1229;
    wire _1230;
    wire _1264;
    wire _1265;
    wire _1266;
    wire _1267;
    wire _1268;
    wire _1269;
    wire _1270;
    wire _1271;
    wire _1272;
    wire _1273;
    wire _1274;
    wire _1275;
    wire _1276;
    wire _1277;
    wire _1278;
    wire _1279;
    wire _1280;
    wire _1281;
    wire _1282;
    wire _1283;
    wire _1284;
    wire _1285;
    wire _1286;
    wire _1287;
    wire _1288;
    wire _1289;
    wire _1290;
    wire _1291;
    wire _1292;
    wire _1293;
    wire _1294;
    wire _1295;
    wire _1329;
    wire _1330;
    wire _1331;
    wire _1332;
    wire _1333;
    wire _1334;
    wire _1335;
    wire _1336;
    wire _1337;
    wire _1338;
    wire _1339;
    wire _1340;
    wire _1341;
    wire _1342;
    wire _1343;
    wire _1344;
    wire _1345;
    wire _1346;
    wire _1347;
    wire _1348;
    wire _1349;
    wire _1350;
    wire _1351;
    wire _1352;
    wire _1353;
    wire _1354;
    wire _1355;
    wire _1356;
    wire _1357;
    wire _1358;
    wire _1359;
    wire _1360;
    wire _1394;
    wire _1395;
    wire _1396;
    wire _1397;
    wire _1398;
    wire _1399;
    wire _1400;
    wire _1401;
    wire _1402;
    wire _1403;
    wire _1404;
    wire _1405;
    wire _1406;
    wire _1407;
    wire _1408;
    wire _1409;
    wire _1410;
    wire _1411;
    wire _1412;
    wire _1413;
    wire _1414;
    wire _1415;
    wire _1416;
    wire _1417;
    wire _1418;
    wire _1419;
    wire _1420;
    wire _1421;
    wire _1422;
    wire _1423;
    wire _1424;
    wire _1425;
    wire _1459;
    wire _1460;
    wire _1461;
    wire _1462;
    wire _1463;
    wire _1464;
    wire _1465;
    wire _1466;
    wire _1467;
    wire _1468;
    wire _1469;
    wire _1470;
    wire _1471;
    wire _1472;
    wire _1473;
    wire _1474;
    wire _1475;
    wire _1476;
    wire _1477;
    wire _1478;
    wire _1479;
    wire _1480;
    wire _1481;
    wire _1482;
    wire _1483;
    wire _1484;
    wire _1485;
    wire _1486;
    wire _1487;
    wire _1488;
    wire _1489;
    wire _1490;
    wire _1524;
    wire _1525;
    wire _1526;
    wire _1527;
    wire _1528;
    wire _1529;
    wire _1530;
    wire _1531;
    wire _1532;
    wire _1533;
    wire _1534;
    wire _1535;
    wire _1536;
    wire _1537;
    wire _1538;
    wire _1539;
    wire _1540;
    wire _1541;
    wire _1542;
    wire _1543;
    wire _1544;
    wire _1545;
    wire _1546;
    wire _1547;
    wire _1548;
    wire _1549;
    wire _1550;
    wire _1551;
    wire _1552;
    wire _1553;
    wire _1554;
    wire _1555;
    wire _1589;
    wire _1590;
    wire _1591;
    wire _1592;
    wire _1593;
    wire _1594;
    wire _1595;
    wire _1596;
    wire _1597;
    wire _1598;
    wire _1599;
    wire _1600;
    wire _1601;
    wire _1602;
    wire _1603;
    wire _1604;
    wire _1605;
    wire _1606;
    wire _1607;
    wire _1608;
    wire _1609;
    wire _1610;
    wire _1611;
    wire _1612;
    wire _1613;
    wire _1614;
    wire _1615;
    wire _1616;
    wire _1617;
    wire _1618;
    wire _1619;
    wire _1620;
    wire _1654;
    wire _1655;
    wire _1656;
    wire _1657;
    wire _1658;
    wire _1659;
    wire _1660;
    wire _1661;
    wire _1662;
    wire _1663;
    wire _1664;
    wire _1665;
    wire _1666;
    wire _1667;
    wire _1668;
    wire _1669;
    wire _1670;
    wire _1671;
    wire _1672;
    wire _1673;
    wire _1674;
    wire _1675;
    wire _1676;
    wire _1677;
    wire _1678;
    wire _1679;
    wire _1680;
    wire _1681;
    wire _1682;
    wire _1683;
    wire _1684;
    wire _1685;
    wire _1719;
    wire _1720;
    wire _1721;
    wire _1722;
    wire _1723;
    wire _1724;
    wire _1725;
    wire _1726;
    wire _1727;
    wire _1728;
    wire _1729;
    wire _1730;
    wire _1731;
    wire _1732;
    wire _1733;
    wire _1734;
    wire _1735;
    wire _1736;
    wire _1737;
    wire _1738;
    wire _1739;
    wire _1740;
    wire _1741;
    wire _1742;
    wire _1743;
    wire _1744;
    wire _1745;
    wire _1746;
    wire _1747;
    wire _1748;
    wire _1749;
    wire _1750;
    wire _1784;
    wire _1785;
    wire _1786;
    wire _1787;
    wire _1788;
    wire _1789;
    wire _1790;
    wire _1791;
    wire _1792;
    wire _1793;
    wire _1794;
    wire _1795;
    wire _1796;
    wire _1797;
    wire _1798;
    wire _1799;
    wire _1800;
    wire _1801;
    wire _1802;
    wire _1803;
    wire _1804;
    wire _1805;
    wire _1806;
    wire _1807;
    wire _1808;
    wire _1809;
    wire _1810;
    wire _1811;
    wire _1812;
    wire _1813;
    wire _1814;
    wire _1815;
    wire _1849;
    wire _1850;
    wire _1851;
    wire _1852;
    wire _1853;
    wire _1854;
    wire _1855;
    wire _1856;
    wire _1857;
    wire _1858;
    wire _1859;
    wire _1860;
    wire _1861;
    wire _1862;
    wire _1863;
    wire _1864;
    wire _1865;
    wire _1866;
    wire _1867;
    wire _1868;
    wire _1869;
    wire _1870;
    wire _1871;
    wire _1872;
    wire _1873;
    wire _1874;
    wire _1875;
    wire _1876;
    wire _1877;
    wire _1878;
    wire _1879;
    wire _1880;
    wire _1914;
    wire _1915;
    wire _1916;
    wire _1917;
    wire _1918;
    wire _1919;
    wire _1920;
    wire _1921;
    wire _1922;
    wire _1923;
    wire _1924;
    wire _1925;
    wire _1926;
    wire _1927;
    wire _1928;
    wire _1929;
    wire _1930;
    wire _1931;
    wire _1932;
    wire _1933;
    wire _1934;
    wire _1935;
    wire _1936;
    wire _1937;
    wire _1938;
    wire _1939;
    wire _1940;
    wire _1941;
    wire _1942;
    wire _1943;
    wire _1944;
    wire _1945;
    wire _1979;
    wire _1980;
    wire _1981;
    wire _1982;
    wire _1983;
    wire _1984;
    wire _1985;
    wire _1986;
    wire _1987;
    wire _1988;
    wire _1989;
    wire _1990;
    wire _1991;
    wire _1992;
    wire _1993;
    wire _1994;
    wire _1995;
    wire _1996;
    wire _1997;
    wire _1998;
    wire _1999;
    wire _2000;
    wire _2001;
    wire _2002;
    wire _2003;
    wire _2004;
    wire _2005;
    wire _2006;
    wire _2007;
    wire _2008;
    wire _2009;
    wire _2010;
    wire _2044;
    wire _2045;
    wire _2046;
    wire _2047;
    wire _2048;
    wire _2049;
    wire _2050;
    wire _2051;
    wire _2052;
    wire _2053;
    wire _2054;
    wire _2055;
    wire _2056;
    wire _2057;
    wire _2058;
    wire _2059;
    wire _2060;
    wire _2061;
    wire _2062;
    wire _2063;
    wire _2064;
    wire _2065;
    wire _2066;
    wire _2067;
    wire _2068;
    wire _2069;
    wire _2070;
    wire _2071;
    wire _2072;
    wire _2073;
    wire _2074;
    wire _2075;
    wire _2109;
    wire _2110;
    wire _2111;
    wire _2112;
    wire _2113;
    wire _2114;
    wire _2115;
    wire _2116;
    wire _2117;
    wire _2118;
    wire _2119;
    wire _2120;
    wire _2121;
    wire _2122;
    wire _2123;
    wire _2124;
    wire _2125;
    wire _2126;
    wire _2127;
    wire _2128;
    wire _2129;
    wire _2130;
    wire _2131;
    wire _2132;
    wire _2133;
    wire _2134;
    wire _2135;
    wire _2136;
    wire _2137;
    wire _2138;
    wire _2139;
    wire _2140;
    wire _2174;
    wire _2175;
    wire _2176;
    wire _2177;
    wire _2178;
    wire _2179;
    wire _2180;
    wire _2181;
    wire _2182;
    wire _2183;
    wire _2184;
    wire _2185;
    wire _2186;
    wire _2187;
    wire _2188;
    wire _2189;
    wire _2190;
    wire _2191;
    wire _2192;
    wire _2193;
    wire _2194;
    wire _2195;
    wire _2196;
    wire _2197;
    wire _2198;
    wire _2199;
    wire _2200;
    wire _2201;
    wire _2202;
    wire _2203;
    wire _2204;
    wire _2205;
    wire _2239;
    wire _2240;
    wire _2241;
    wire _2242;
    wire _2243;
    wire _2244;
    wire _2245;
    wire _2246;
    wire _2247;
    wire _2248;
    wire _2249;
    wire _2250;
    wire _2251;
    wire _2252;
    wire _2253;
    wire _2254;
    wire _2255;
    wire _2256;
    wire _2257;
    wire _2258;
    wire _2259;
    wire _2260;
    wire _2261;
    wire _2262;
    wire _2263;
    wire _2264;
    wire _2265;
    wire _2266;
    wire _2267;
    wire _2268;
    wire _2269;
    wire _2270;
    wire _2304;
    wire _2305;
    wire _2306;
    wire _2307;
    wire _2308;
    wire _2309;
    wire _2310;
    wire _2311;
    wire _2312;
    wire _2313;
    wire _2314;
    wire _2315;
    wire _2316;
    wire _2317;
    wire _2318;
    wire _2319;
    wire _2320;
    wire _2321;
    wire _2322;
    wire _2323;
    wire _2324;
    wire _2325;
    wire _2326;
    wire _2327;
    wire _2328;
    wire _2329;
    wire _2330;
    wire _2331;
    wire _2332;
    wire _2333;
    wire _2334;
    wire _2335;
    wire _2369;
    wire _2370;
    wire _2371;
    wire _2372;
    wire _2373;
    wire _2374;
    wire _2375;
    wire _2376;
    wire _2377;
    wire _2378;
    wire _2379;
    wire _2380;
    wire _2381;
    wire _2382;
    wire _2383;
    wire _2384;
    wire _2385;
    wire _2386;
    wire _2387;
    wire _2388;
    wire _2389;
    wire _2390;
    wire _2391;
    wire _2392;
    wire _2393;
    wire _2394;
    wire _2395;
    wire _2396;
    wire _2397;
    wire _2398;
    wire _2399;
    wire _2400;
    wire _2434;
    wire _2435;
    wire _2436;
    wire _2437;
    wire _2438;
    wire _2439;
    wire _2440;
    wire _2441;
    wire _2442;
    wire _2443;
    wire _2444;
    wire _2445;
    wire _2446;
    wire _2447;
    wire _2448;
    wire _2449;
    wire _2450;
    wire _2451;
    wire _2452;
    wire _2453;
    wire _2454;
    wire _2455;
    wire _2456;
    wire _2457;
    wire _2458;
    wire _2459;
    wire _2460;
    wire _2461;
    wire _2462;
    wire _2463;
    wire _2464;
    wire _2465;
    wire _2499;
    wire _2500;
    wire _2501;
    wire _2502;
    wire _2503;
    wire _2504;
    wire _2505;
    wire _2506;
    wire _2507;
    wire _2508;
    wire _2509;
    wire _2510;
    wire _2511;
    wire _2512;
    wire _2513;
    wire _2514;
    wire _2515;
    wire _2516;
    wire _2517;
    wire _2518;
    wire _2519;
    wire _2520;
    wire _2521;
    wire _2522;
    wire _2523;
    wire _2524;
    wire _2525;
    wire _2526;
    wire _2527;
    wire _2528;
    wire _2529;
    wire _2530;
    wire _2564;
    wire _2565;
    wire _2566;
    wire _2567;
    wire _2568;
    wire _2569;
    wire _2570;
    wire _2571;
    wire _2572;
    wire _2573;
    wire _2574;
    wire _2575;
    wire _2576;
    wire _2577;
    wire _2578;
    wire _2579;
    wire _2580;
    wire _2581;
    wire _2582;
    wire _2583;
    wire _2584;
    wire _2585;
    wire _2586;
    wire _2587;
    wire _2588;
    wire _2589;
    wire _2590;
    wire _2591;
    wire _2592;
    wire _2593;
    wire _2594;
    wire _2595;
    wire _2629;
    wire _2630;
    wire _2631;
    wire _2632;
    wire _2633;
    wire _2634;
    wire _2635;
    wire _2636;
    wire _2637;
    wire _2638;
    wire _2639;
    wire _2640;
    wire _2641;
    wire _2642;
    wire _2643;
    wire _2644;
    wire _2645;
    wire _2646;
    wire _2647;
    wire _2648;
    wire _2649;
    wire _2650;
    wire _2651;
    wire _2652;
    wire _2653;
    wire _2654;
    wire _2655;
    wire _2656;
    wire _2657;
    wire _2658;
    wire _2659;
    wire _2660;
    wire _2694;
    wire _2695;
    wire _2696;
    wire _2697;
    wire _2698;
    wire _2699;
    wire _2700;
    wire _2701;
    wire _2702;
    wire _2703;
    wire _2704;
    wire _2705;
    wire _2706;
    wire _2707;
    wire _2708;
    wire _2709;
    wire _2710;
    wire _2711;
    wire _2712;
    wire _2713;
    wire _2714;
    wire _2715;
    wire _2716;
    wire _2717;
    wire _2718;
    wire _2719;
    wire _2720;
    wire _2721;
    wire _2722;
    wire _2723;
    wire _2724;
    wire _2725;
    wire _2759;
    wire _2760;
    wire _2761;
    wire _2762;
    wire _2763;
    wire _2764;
    wire _2765;
    wire _2766;
    wire _2767;
    wire _2768;
    wire _2769;
    wire _2770;
    wire _2771;
    wire _2772;
    wire _2773;
    wire _2774;
    wire _2775;
    wire _2776;
    wire _2777;
    wire _2778;
    wire _2779;
    wire _2780;
    wire _2781;
    wire _2782;
    wire _2783;
    wire _2784;
    wire _2785;
    wire _2786;
    wire _2787;
    wire _2788;
    wire _2789;
    wire _2790;
    wire _2824;
    wire _2825;
    wire _2826;
    wire _2827;
    wire _2828;
    wire _2829;
    wire _2830;
    wire _2831;
    wire _2832;
    wire _2833;
    wire _2834;
    wire _2835;
    wire _2836;
    wire _2837;
    wire _2838;
    wire _2839;
    wire _2840;
    wire _2841;
    wire _2842;
    wire _2843;
    wire _2844;
    wire _2845;
    wire _2846;
    wire _2847;
    wire _2848;
    wire _2849;
    wire _2850;
    wire _2851;
    wire _2852;
    wire _2853;
    wire _2854;
    wire _2855;
    wire _2889;
    wire _2890;
    wire _2891;
    wire _2892;
    wire _2893;
    wire _2894;
    wire _2895;
    wire _2896;
    wire _2897;
    wire _2898;
    wire _2899;
    wire _2900;
    wire _2901;
    wire _2902;
    wire _2903;
    wire _2904;
    wire _2905;
    wire _2906;
    wire _2907;
    wire _2908;
    wire _2909;
    wire _2910;
    wire _2911;
    wire _2912;
    wire _2913;
    wire _2914;
    wire _2915;
    wire _2916;
    wire _2917;
    wire _2918;
    wire _2919;
    wire _2920;
    wire _2954;
    wire _2955;
    wire _2956;
    wire _2957;
    wire _2958;
    wire _2959;
    wire _2960;
    wire _2961;
    wire _2962;
    wire _2963;
    wire _2964;
    wire _2965;
    wire _2966;
    wire _2967;
    wire _2968;
    wire _2969;
    wire _2970;
    wire _2971;
    wire _2972;
    wire _2973;
    wire _2974;
    wire _2975;
    wire _2976;
    wire _2977;
    wire _2978;
    wire _2979;
    wire _2980;
    wire _2981;
    wire _2982;
    wire _2983;
    wire _2984;
    wire _2985;
    wire _3019;
    wire _3020;
    wire _3021;
    wire _3022;
    wire _3023;
    wire _3024;
    wire _3025;
    wire _3026;
    wire _3027;
    wire _3028;
    wire _3029;
    wire _3030;
    wire _3031;
    wire _3032;
    wire _3033;
    wire _3034;
    wire _3035;
    wire _3036;
    wire _3037;
    wire _3038;
    wire _3039;
    wire _3040;
    wire _3041;
    wire _3042;
    wire _3043;
    wire _3044;
    wire _3045;
    wire _3046;
    wire _3047;
    wire _3048;
    wire _3049;
    wire _3050;
    wire _3084;
    wire _3085;
    wire _3086;
    wire _3087;
    wire _3088;
    wire _3089;
    wire _3090;
    wire _3091;
    wire _3092;
    wire _3093;
    wire _3094;
    wire _3095;
    wire _3096;
    wire _3097;
    wire _3098;
    wire _3099;
    wire _3100;
    wire _3101;
    wire _3102;
    wire _3103;
    wire _3104;
    wire _3105;
    wire _3106;
    wire _3107;
    wire _3108;
    wire _3109;
    wire _3110;
    wire _3111;
    wire _3112;
    wire _3113;
    wire _3114;
    wire _3115;
    wire _3149;
    wire _3150;
    wire _3151;
    wire _3152;
    wire _3153;
    wire _3154;
    wire _3155;
    wire _3156;
    wire _3157;
    wire _3158;
    wire _3159;
    wire _3160;
    wire _3161;
    wire _3162;
    wire _3163;
    wire _3164;
    wire _3165;
    wire _3166;
    wire _3167;
    wire _3168;
    wire _3169;
    wire _3170;
    wire _3171;
    wire _3172;
    wire _3173;
    wire _3174;
    wire _3175;
    wire _3176;
    wire _3177;
    wire _3178;
    wire _3179;
    wire _3180;
    wire _3214;
    wire _3215;
    wire _3216;
    wire _3217;
    wire _3218;
    wire _3219;
    wire _3220;
    wire _3221;
    wire _3222;
    wire _3223;
    wire _3224;
    wire _3225;
    wire _3226;
    wire _3227;
    wire _3228;
    wire _3229;
    wire _3230;
    wire _3231;
    wire _3232;
    wire _3233;
    wire _3234;
    wire _3235;
    wire _3236;
    wire _3237;
    wire _3238;
    wire _3239;
    wire _3240;
    wire _3241;
    wire _3242;
    wire _3243;
    wire _3244;
    wire _3245;
    wire _3279;
    wire _3280;
    wire _3281;
    wire _3282;
    wire _3283;
    wire _3284;
    wire _3285;
    wire _3286;
    wire _3287;
    wire _3288;
    wire _3289;
    wire _3290;
    wire _3291;
    wire _3292;
    wire _3293;
    wire _3294;
    wire _3295;
    wire _3296;
    wire _3297;
    wire _3298;
    wire _3299;
    wire _3300;
    wire _3301;
    wire _3302;
    wire _3303;
    wire _3304;
    wire _3305;
    wire _3306;
    wire _3307;
    wire _3308;
    wire _3309;
    wire _3310;
    wire _3344;
    wire _3345;
    wire _3346;
    wire _3347;
    wire _3348;
    wire _3349;
    wire _3350;
    wire _3351;
    wire _3352;
    wire _3353;
    wire _3354;
    wire _3355;
    wire _3356;
    wire _3357;
    wire _3358;
    wire _3359;
    wire _3360;
    wire _3361;
    wire _3362;
    wire _3363;
    wire _3364;
    wire _3365;
    wire _3366;
    wire _3367;
    wire _3368;
    wire _3369;
    wire _3370;
    wire _3371;
    wire _3372;
    wire _3373;
    wire _3374;
    wire _3375;
    wire _3409;
    wire _3410;
    wire _3411;
    wire _3412;
    wire _3413;
    wire _3414;
    wire _3415;
    wire _3416;
    wire _3417;
    wire _3418;
    wire _3419;
    wire _3420;
    wire _3421;
    wire _3422;
    wire _3423;
    wire _3424;
    wire _3425;
    wire _3426;
    wire _3427;
    wire _3428;
    wire _3429;
    wire _3430;
    wire _3431;
    wire _3432;
    wire _3433;
    wire _3434;
    wire _3435;
    wire _3436;
    wire _3437;
    wire _3438;
    wire _3439;
    wire _3440;
    wire _3474;
    wire _3475;
    wire _3476;
    wire _3477;
    wire _3478;
    wire _3479;
    wire _3480;
    wire _3481;
    wire _3482;
    wire _3483;
    wire _3484;
    wire _3485;
    wire _3486;
    wire _3487;
    wire _3488;
    wire _3489;
    wire _3490;
    wire _3491;
    wire _3492;
    wire _3493;
    wire _3494;
    wire _3495;
    wire _3496;
    wire _3497;
    wire _3498;
    wire _3499;
    wire _3500;
    wire _3501;
    wire _3502;
    wire _3503;
    wire _3504;
    wire _3505;
    wire _3539;
    wire _3540;
    wire _3541;
    wire _3542;
    wire _3543;
    wire _3544;
    wire _3545;
    wire _3546;
    wire _3547;
    wire _3548;
    wire _3549;
    wire _3550;
    wire _3551;
    wire _3552;
    wire _3553;
    wire _3554;
    wire _3555;
    wire _3556;
    wire _3557;
    wire _3558;
    wire _3559;
    wire _3560;
    wire _3561;
    wire _3562;
    wire _3563;
    wire _3564;
    wire _3565;
    wire _3566;
    wire _3567;
    wire _3568;
    wire _3569;
    wire _3570;
    wire _3604;
    wire _3605;
    wire _3606;
    wire _3607;
    wire _3608;
    wire _3609;
    wire _3610;
    wire _3611;
    wire _3612;
    wire _3613;
    wire _3614;
    wire _3615;
    wire _3616;
    wire _3617;
    wire _3618;
    wire _3619;
    wire _3620;
    wire _3621;
    wire _3622;
    wire _3623;
    wire _3624;
    wire _3625;
    wire _3626;
    wire _3627;
    wire _3628;
    wire _3629;
    wire _3630;
    wire _3631;
    wire _3632;
    wire _3633;
    wire _3634;
    wire _3635;
    wire _3669;
    wire _3670;
    wire _3671;
    wire _3672;
    wire _3673;
    wire _3674;
    wire _3675;
    wire _3676;
    wire _3677;
    wire _3678;
    wire _3679;
    wire _3680;
    wire _3681;
    wire _3682;
    wire _3683;
    wire _3684;
    wire _3685;
    wire _3686;
    wire _3687;
    wire _3688;
    wire _3689;
    wire _3690;
    wire _3691;
    wire _3692;
    wire _3693;
    wire _3694;
    wire _3695;
    wire _3696;
    wire _3697;
    wire _3698;
    wire _3699;
    wire _3700;
    wire _3734;
    wire _3735;
    wire _3736;
    wire _3737;
    wire _3738;
    wire _3739;
    wire _3740;
    wire _3741;
    wire _3742;
    wire _3743;
    wire _3744;
    wire _3745;
    wire _3746;
    wire _3747;
    wire _3748;
    wire _3749;
    wire _3750;
    wire _3751;
    wire _3752;
    wire _3753;
    wire _3754;
    wire _3755;
    wire _3756;
    wire _3757;
    wire _3758;
    wire _3759;
    wire _3760;
    wire _3761;
    wire _3762;
    wire _3763;
    wire _3764;
    wire _3765;
    wire _3799;
    wire _3800;
    wire _3801;
    wire _3802;
    wire _3803;
    wire _3804;
    wire _3805;
    wire _3806;
    wire _3807;
    wire _3808;
    wire _3809;
    wire _3810;
    wire _3811;
    wire _3812;
    wire _3813;
    wire _3814;
    wire _3815;
    wire _3816;
    wire _3817;
    wire _3818;
    wire _3819;
    wire _3820;
    wire _3821;
    wire _3822;
    wire _3823;
    wire _3824;
    wire _3825;
    wire _3826;
    wire _3827;
    wire _3828;
    wire _3829;
    wire _3830;
    wire _3864;
    wire _3865;
    wire _3866;
    wire _3867;
    wire _3868;
    wire _3869;
    wire _3870;
    wire _3871;
    wire _3872;
    wire _3873;
    wire _3874;
    wire _3875;
    wire _3876;
    wire _3877;
    wire _3878;
    wire _3879;
    wire _3880;
    wire _3881;
    wire _3882;
    wire _3883;
    wire _3884;
    wire _3885;
    wire _3886;
    wire _3887;
    wire _3888;
    wire _3889;
    wire _3890;
    wire _3891;
    wire _3892;
    wire _3893;
    wire _3894;
    wire _3895;
    wire _3929;
    wire _3930;
    wire _3931;
    wire _3932;
    wire _3933;
    wire _3934;
    wire _3935;
    wire _3936;
    wire _3937;
    wire _3938;
    wire _3939;
    wire _3940;
    wire _3941;
    wire _3942;
    wire _3943;
    wire _3944;
    wire _3945;
    wire _3946;
    wire _3947;
    wire _3948;
    wire _3949;
    wire _3950;
    wire _3951;
    wire _3952;
    wire _3953;
    wire _3954;
    wire _3955;
    wire _3956;
    wire _3957;
    wire _3958;
    wire _3959;
    wire _3960;
    wire _3994;
    wire _3995;
    wire _3996;
    wire _3997;
    wire _3998;
    wire _3999;
    wire _4000;
    wire _4001;
    wire _4002;
    wire _4003;
    wire _4004;
    wire _4005;
    wire _4006;
    wire _4007;
    wire _4008;
    wire _4009;
    wire _4010;
    wire _4011;
    wire _4012;
    wire _4013;
    wire _4014;
    wire _4015;
    wire _4016;
    wire _4017;
    wire _4018;
    wire _4019;
    wire _4020;
    wire _4021;
    wire _4022;
    wire _4023;
    wire _4024;
    wire _4025;
    wire _4059;
    wire _4060;
    wire _4061;
    wire _4062;
    wire _4063;
    wire _4064;
    wire _4065;
    wire _4066;
    wire _4067;
    wire _4068;
    wire _4069;
    wire _4070;
    wire _4071;
    wire _4072;
    wire _4073;
    wire _4074;
    wire _4075;
    wire _4076;
    wire _4077;
    wire _4078;
    wire _4079;
    wire _4080;
    wire _4081;
    wire _4082;
    wire _4083;
    wire _4084;
    wire _4085;
    wire _4086;
    wire _4087;
    wire _4088;
    wire _4089;
    wire _4090;
    wire _4124;
    wire _4125;
    wire _4126;
    wire _4127;
    wire _4128;
    wire _4129;
    wire _4130;
    wire _4131;
    wire _4132;
    wire _4133;
    wire _4134;
    wire _4135;
    wire _4136;
    wire _4137;
    wire _4138;
    wire _4139;
    wire _4140;
    wire _4141;
    wire _4142;
    wire _4143;
    wire _4144;
    wire _4145;
    wire _4146;
    wire _4147;
    wire _4148;
    wire _4149;
    wire _4150;
    wire _4151;
    wire _4152;
    wire _4153;
    wire _4154;
    wire _4155;
    wire _4189;
    wire _4190;
    wire _4191;
    wire _4192;
    wire _4193;
    wire _4194;
    wire _4195;
    wire _4196;
    wire _4197;
    wire _4198;
    wire _4199;
    wire _4200;
    wire _4201;
    wire _4202;
    wire _4203;
    wire _4204;
    wire _4205;
    wire _4206;
    wire _4207;
    wire _4208;
    wire _4209;
    wire _4210;
    wire _4211;
    wire _4212;
    wire _4213;
    wire _4214;
    wire _4215;
    wire _4216;
    wire _4217;
    wire _4218;
    wire _4219;
    wire _4220;
    wire _4254;
    wire _4255;
    wire _4256;
    wire _4257;
    wire _4258;
    wire _4259;
    wire _4260;
    wire _4261;
    wire _4262;
    wire _4263;
    wire _4264;
    wire _4265;
    wire _4266;
    wire _4267;
    wire _4268;
    wire _4269;
    wire _4270;
    wire _4271;
    wire _4272;
    wire _4273;
    wire _4274;
    wire _4275;
    wire _4276;
    wire _4277;
    wire _4278;
    wire _4279;
    wire _4280;
    wire _4281;
    wire _4282;
    wire _4283;
    wire _4284;
    wire _4285;
    wire _4319;
    wire _4320;
    wire _4321;
    wire _4322;
    wire _4323;
    wire _4324;
    wire _4325;
    wire _4326;
    wire _4327;
    wire _4328;
    wire _4329;
    wire _4330;
    wire _4331;
    wire _4332;
    wire _4333;
    wire _4334;
    wire _4335;
    wire _4336;
    wire _4337;
    wire _4338;
    wire _4339;
    wire _4340;
    wire _4341;
    wire _4342;
    wire _4343;
    wire _4344;
    wire _4345;
    wire _4346;
    wire _4347;
    wire _4348;
    wire _4349;
    wire _4350;
    wire _4384;
    wire _4385;
    wire _4386;
    wire _4387;
    wire _4388;
    wire _4389;
    wire _4390;
    wire _4391;
    wire _4392;
    wire _4393;
    wire _4394;
    wire _4395;
    wire _4396;
    wire _4397;
    wire _4398;
    wire _4399;
    wire _4400;
    wire _4401;
    wire _4402;
    wire _4403;
    wire _4404;
    wire _4405;
    wire _4406;
    wire _4407;
    wire _4408;
    wire _4409;
    wire _4410;
    wire _4411;
    wire _4412;
    wire _4413;
    wire _4414;
    wire _4415;
    wire _4449;
    wire _4450;
    wire _4451;
    wire _4452;
    wire _4453;
    wire _4454;
    wire _4455;
    wire _4456;
    wire _4457;
    wire _4458;
    wire _4459;
    wire _4460;
    wire _4461;
    wire _4462;
    wire _4463;
    wire _4464;
    wire _4465;
    wire _4466;
    wire _4467;
    wire _4468;
    wire _4469;
    wire _4470;
    wire _4471;
    wire _4472;
    wire _4473;
    wire _4474;
    wire _4475;
    wire _4476;
    wire _4477;
    wire _4478;
    wire _4479;
    wire _4480;
    wire _4514;
    wire _4515;
    wire _4516;
    wire _4517;
    wire _4518;
    wire _4519;
    wire _4520;
    wire _4521;
    wire _4522;
    wire _4523;
    wire _4524;
    wire _4525;
    wire _4526;
    wire _4527;
    wire _4528;
    wire _4529;
    wire _4530;
    wire _4531;
    wire _4532;
    wire _4533;
    wire _4534;
    wire _4535;
    wire _4536;
    wire _4537;
    wire _4538;
    wire _4539;
    wire _4540;
    wire _4541;
    wire _4542;
    wire _4543;
    wire _4544;
    wire _4545;
    wire _4579;
    wire _4580;
    wire _4581;
    wire _4582;
    wire _4583;
    wire _4584;
    wire _4585;
    wire _4586;
    wire _4587;
    wire _4588;
    wire _4589;
    wire _4590;
    wire _4591;
    wire _4592;
    wire _4593;
    wire _4594;
    wire _4595;
    wire _4596;
    wire _4597;
    wire _4598;
    wire _4599;
    wire _4600;
    wire _4601;
    wire _4602;
    wire _4603;
    wire _4604;
    wire _4605;
    wire _4606;
    wire _4607;
    wire _4608;
    wire _4609;
    wire _4610;
    wire _4644;
    wire _4645;
    wire _4646;
    wire _4647;
    wire _4648;
    wire _4649;
    wire _4650;
    wire _4651;
    wire _4652;
    wire _4653;
    wire _4654;
    wire _4655;
    wire _4656;
    wire _4657;
    wire _4658;
    wire _4659;
    wire _4660;
    wire _4661;
    wire _4662;
    wire _4663;
    wire _4664;
    wire _4665;
    wire _4666;
    wire _4667;
    wire _4668;
    wire _4669;
    wire _4670;
    wire _4671;
    wire _4672;
    wire _4673;
    wire _4674;
    wire _4675;
    wire _4709;
    wire _4710;
    wire _4711;
    wire _4712;
    wire _4713;
    wire _4714;
    wire _4715;
    wire _4716;
    wire _4717;
    wire _4718;
    wire _4719;
    wire _4720;
    wire _4721;
    wire _4722;
    wire _4723;
    wire _4724;
    wire _4725;
    wire _4726;
    wire _4727;
    wire _4728;
    wire _4729;
    wire _4730;
    wire _4731;
    wire _4732;
    wire _4733;
    wire _4734;
    wire _4735;
    wire _4736;
    wire _4737;
    wire _4738;
    wire _4739;
    wire _4740;
    wire _4774;
    wire _4775;
    wire _4776;
    wire _4777;
    wire _4778;
    wire _4779;
    wire _4780;
    wire _4781;
    wire _4782;
    wire _4783;
    wire _4784;
    wire _4785;
    wire _4786;
    wire _4787;
    wire _4788;
    wire _4789;
    wire _4790;
    wire _4791;
    wire _4792;
    wire _4793;
    wire _4794;
    wire _4795;
    wire _4796;
    wire _4797;
    wire _4798;
    wire _4799;
    wire _4800;
    wire _4801;
    wire _4802;
    wire _4803;
    wire _4804;
    wire _4805;
    wire _4839;
    wire _4840;
    wire _4841;
    wire _4842;
    wire _4843;
    wire _4844;
    wire _4845;
    wire _4846;
    wire _4847;
    wire _4848;
    wire _4849;
    wire _4850;
    wire _4851;
    wire _4852;
    wire _4853;
    wire _4854;
    wire _4855;
    wire _4856;
    wire _4857;
    wire _4858;
    wire _4859;
    wire _4860;
    wire _4861;
    wire _4862;
    wire _4863;
    wire _4864;
    wire _4865;
    wire _4866;
    wire _4867;
    wire _4868;
    wire _4869;
    wire _4870;
    wire _4904;
    wire _4905;
    wire _4906;
    wire _4907;
    wire _4908;
    wire _4909;
    wire _4910;
    wire _4911;
    wire _4912;
    wire _4913;
    wire _4914;
    wire _4915;
    wire _4916;
    wire _4917;
    wire _4918;
    wire _4919;
    wire _4920;
    wire _4921;
    wire _4922;
    wire _4923;
    wire _4924;
    wire _4925;
    wire _4926;
    wire _4927;
    wire _4928;
    wire _4929;
    wire _4930;
    wire _4931;
    wire _4932;
    wire _4933;
    wire _4934;
    wire _4935;
    wire _4969;
    wire _4970;
    wire _4971;
    wire _4972;
    wire _4973;
    wire _4974;
    wire _4975;
    wire _4976;
    wire _4977;
    wire _4978;
    wire _4979;
    wire _4980;
    wire _4981;
    wire _4982;
    wire _4983;
    wire _4984;
    wire _4985;
    wire _4986;
    wire _4987;
    wire _4988;
    wire _4989;
    wire _4990;
    wire _4991;
    wire _4992;
    wire _4993;
    wire _4994;
    wire _4995;
    wire _4996;
    wire _4997;
    wire _4998;
    wire _4999;
    wire _5000;
    wire _5034;
    wire _5035;
    wire _5036;
    wire _5037;
    wire _5038;
    wire _5039;
    wire _5040;
    wire _5041;
    wire _5042;
    wire _5043;
    wire _5044;
    wire _5045;
    wire _5046;
    wire _5047;
    wire _5048;
    wire _5049;
    wire _5050;
    wire _5051;
    wire _5052;
    wire _5053;
    wire _5054;
    wire _5055;
    wire _5056;
    wire _5057;
    wire _5058;
    wire _5059;
    wire _5060;
    wire _5061;
    wire _5062;
    wire _5063;
    wire _5064;
    wire _5065;
    wire _5099;
    wire _5100;
    wire _5101;
    wire _5102;
    wire _5103;
    wire _5104;
    wire _5105;
    wire _5106;
    wire _5107;
    wire _5108;
    wire _5109;
    wire _5110;
    wire _5111;
    wire _5112;
    wire _5113;
    wire _5114;
    wire _5115;
    wire _5116;
    wire _5117;
    wire _5118;
    wire _5119;
    wire _5120;
    wire _5121;
    wire _5122;
    wire _5123;
    wire _5124;
    wire _5125;
    wire _5126;
    wire _5127;
    wire _5128;
    wire _5129;
    wire _5130;
    wire _5164;
    wire _5165;
    wire _5166;
    wire _5167;
    wire _5168;
    wire _5169;
    wire _5170;
    wire _5171;
    wire _5172;
    wire _5173;
    wire _5174;
    wire _5175;
    wire _5176;
    wire _5177;
    wire _5178;
    wire _5179;
    wire _5180;
    wire _5181;
    wire _5182;
    wire _5183;
    wire _5184;
    wire _5185;
    wire _5186;
    wire _5187;
    wire _5188;
    wire _5189;
    wire _5190;
    wire _5191;
    wire _5192;
    wire _5193;
    wire _5194;
    wire _5195;
    wire _5229;
    wire _5230;
    wire _5231;
    wire _5232;
    wire _5233;
    wire _5234;
    wire _5235;
    wire _5236;
    wire _5237;
    wire _5238;
    wire _5239;
    wire _5240;
    wire _5241;
    wire _5242;
    wire _5243;
    wire _5244;
    wire _5245;
    wire _5246;
    wire _5247;
    wire _5248;
    wire _5249;
    wire _5250;
    wire _5251;
    wire _5252;
    wire _5253;
    wire _5254;
    wire _5255;
    wire _5256;
    wire _5257;
    wire _5258;
    wire _5259;
    wire _5260;
    wire _5294;
    wire _5295;
    wire _5296;
    wire _5297;
    wire _5298;
    wire _5299;
    wire _5300;
    wire _5301;
    wire _5302;
    wire _5303;
    wire _5304;
    wire _5305;
    wire _5306;
    wire _5307;
    wire _5308;
    wire _5309;
    wire _5310;
    wire _5311;
    wire _5312;
    wire _5313;
    wire _5314;
    wire _5315;
    wire _5316;
    wire _5317;
    wire _5318;
    wire _5319;
    wire _5320;
    wire _5321;
    wire _5322;
    wire _5323;
    wire _5324;
    wire _5325;
    wire _5359;
    wire _5360;
    wire _5361;
    wire _5362;
    wire _5363;
    wire _5364;
    wire _5365;
    wire _5366;
    wire _5367;
    wire _5368;
    wire _5369;
    wire _5370;
    wire _5371;
    wire _5372;
    wire _5373;
    wire _5374;
    wire _5375;
    wire _5376;
    wire _5377;
    wire _5378;
    wire _5379;
    wire _5380;
    wire _5381;
    wire _5382;
    wire _5383;
    wire _5384;
    wire _5385;
    wire _5386;
    wire _5387;
    wire _5388;
    wire _5389;
    wire _5390;
    wire _5424;
    wire _5425;
    wire _5426;
    wire _5427;
    wire _5428;
    wire _5429;
    wire _5430;
    wire _5431;
    wire _5432;
    wire _5433;
    wire _5434;
    wire _5435;
    wire _5436;
    wire _5437;
    wire _5438;
    wire _5439;
    wire _5440;
    wire _5441;
    wire _5442;
    wire _5443;
    wire _5444;
    wire _5445;
    wire _5446;
    wire _5447;
    wire _5448;
    wire _5449;
    wire _5450;
    wire _5451;
    wire _5452;
    wire _5453;
    wire _5454;
    wire _5455;
    assign _0 = \a[0][0] ;
    assign _1 = \a[0][1] ;
    assign _2 = \a[0][2] ;
    assign _3 = \a[0][3] ;
    assign _4 = \a[0][4] ;
    assign _5 = \a[0][5] ;
    assign _6 = \a[0][6] ;
    assign _7 = \a[0][7] ;
    assign _8 = \a[0][8] ;
    assign _9 = \a[0][9] ;
    assign _10 = \a[0][10] ;
    assign _11 = \a[0][11] ;
    assign _12 = \a[0][12] ;
    assign _13 = \a[0][13] ;
    assign _14 = \a[0][14] ;
    assign _15 = \a[0][15] ;
    assign _16 = \a[1][0] ;
    assign _17 = \a[1][1] ;
    assign _18 = \a[1][2] ;
    assign _19 = \a[1][3] ;
    assign _20 = \a[1][4] ;
    assign _21 = \a[1][5] ;
    assign _22 = \a[1][6] ;
    assign _23 = \a[1][7] ;
    assign _24 = \a[1][8] ;
    assign _25 = \a[1][9] ;
    assign _26 = \a[1][10] ;
    assign _27 = \a[1][11] ;
    assign _28 = \a[1][12] ;
    assign _29 = \a[1][13] ;
    assign _30 = \a[1][14] ;
    assign _31 = \a[1][15] ;
    assign _32 = \a[2][0] ;
    assign _33 = \a[2][1] ;
    assign _34 = \a[2][2] ;
    assign _35 = \a[2][3] ;
    assign _36 = \a[2][4] ;
    assign _37 = \a[2][5] ;
    assign _38 = \a[2][6] ;
    assign _39 = \a[2][7] ;
    assign _40 = \a[2][8] ;
    assign _41 = \a[2][9] ;
    assign _42 = \a[2][10] ;
    assign _43 = \a[2][11] ;
    assign _44 = \a[2][12] ;
    assign _45 = \a[2][13] ;
    assign _46 = \a[2][14] ;
    assign _47 = \a[2][15] ;
    assign _48 = \a[3][0] ;
    assign _49 = \a[3][1] ;
    assign _50 = \a[3][2] ;
    assign _51 = \a[3][3] ;
    assign _52 = \a[3][4] ;
    assign _53 = \a[3][5] ;
    assign _54 = \a[3][6] ;
    assign _55 = \a[3][7] ;
    assign _56 = \a[3][8] ;
    assign _57 = \a[3][9] ;
    assign _58 = \a[3][10] ;
    assign _59 = \a[3][11] ;
    assign _60 = \a[3][12] ;
    assign _61 = \a[3][13] ;
    assign _62 = \a[3][14] ;
    assign _63 = \a[3][15] ;
    assign _64 = \a[4][0] ;
    assign _65 = \a[4][1] ;
    assign _66 = \a[4][2] ;
    assign _67 = \a[4][3] ;
    assign _68 = \a[4][4] ;
    assign _69 = \a[4][5] ;
    assign _70 = \a[4][6] ;
    assign _71 = \a[4][7] ;
    assign _72 = \a[4][8] ;
    assign _73 = \a[4][9] ;
    assign _74 = \a[4][10] ;
    assign _75 = \a[4][11] ;
    assign _76 = \a[4][12] ;
    assign _77 = \a[4][13] ;
    assign _78 = \a[4][14] ;
    assign _79 = \a[4][15] ;
    assign _80 = \a[5][0] ;
    assign _81 = \a[5][1] ;
    assign _82 = \a[5][2] ;
    assign _83 = \a[5][3] ;
    assign _84 = \a[5][4] ;
    assign _85 = \a[5][5] ;
    assign _86 = \a[5][6] ;
    assign _87 = \a[5][7] ;
    assign _88 = \a[5][8] ;
    assign _89 = \a[5][9] ;
    assign _90 = \a[5][10] ;
    assign _91 = \a[5][11] ;
    assign _92 = \a[5][12] ;
    assign _93 = \a[5][13] ;
    assign _94 = \a[5][14] ;
    assign _95 = \a[5][15] ;
    assign _96 = \a[6][0] ;
    assign _97 = \a[6][1] ;
    assign _98 = \a[6][2] ;
    assign _99 = \a[6][3] ;
    assign _100 = \a[6][4] ;
    assign _101 = \a[6][5] ;
    assign _102 = \a[6][6] ;
    assign _103 = \a[6][7] ;
    assign _104 = \a[6][8] ;
    assign _105 = \a[6][9] ;
    assign _106 = \a[6][10] ;
    assign _107 = \a[6][11] ;
    assign _108 = \a[6][12] ;
    assign _109 = \a[6][13] ;
    assign _110 = \a[6][14] ;
    assign _111 = \a[6][15] ;
    assign _112 = \a[7][0] ;
    assign _113 = \a[7][1] ;
    assign _114 = \a[7][2] ;
    assign _115 = \a[7][3] ;
    assign _116 = \a[7][4] ;
    assign _117 = \a[7][5] ;
    assign _118 = \a[7][6] ;
    assign _119 = \a[7][7] ;
    assign _120 = \a[7][8] ;
    assign _121 = \a[7][9] ;
    assign _122 = \a[7][10] ;
    assign _123 = \a[7][11] ;
    assign _124 = \a[7][12] ;
    assign _125 = \a[7][13] ;
    assign _126 = \a[7][14] ;
    assign _127 = \a[7][15] ;
    assign _128 = \a[8][0] ;
    assign _129 = \a[8][1] ;
    assign _130 = \a[8][2] ;
    assign _131 = \a[8][3] ;
    assign _132 = \a[8][4] ;
    assign _133 = \a[8][5] ;
    assign _134 = \a[8][6] ;
    assign _135 = \a[8][7] ;
    assign _136 = \a[8][8] ;
    assign _137 = \a[8][9] ;
    assign _138 = \a[8][10] ;
    assign _139 = \a[8][11] ;
    assign _140 = \a[8][12] ;
    assign _141 = \a[8][13] ;
    assign _142 = \a[8][14] ;
    assign _143 = \a[8][15] ;
    assign _144 = \a[9][0] ;
    assign _145 = \a[9][1] ;
    assign _146 = \a[9][2] ;
    assign _147 = \a[9][3] ;
    assign _148 = \a[9][4] ;
    assign _149 = \a[9][5] ;
    assign _150 = \a[9][6] ;
    assign _151 = \a[9][7] ;
    assign _152 = \a[9][8] ;
    assign _153 = \a[9][9] ;
    assign _154 = \a[9][10] ;
    assign _155 = \a[9][11] ;
    assign _156 = \a[9][12] ;
    assign _157 = \a[9][13] ;
    assign _158 = \a[9][14] ;
    assign _159 = \a[9][15] ;
    assign _160 = \a[10][0] ;
    assign _161 = \a[10][1] ;
    assign _162 = \a[10][2] ;
    assign _163 = \a[10][3] ;
    assign _164 = \a[10][4] ;
    assign _165 = \a[10][5] ;
    assign _166 = \a[10][6] ;
    assign _167 = \a[10][7] ;
    assign _168 = \a[10][8] ;
    assign _169 = \a[10][9] ;
    assign _170 = \a[10][10] ;
    assign _171 = \a[10][11] ;
    assign _172 = \a[10][12] ;
    assign _173 = \a[10][13] ;
    assign _174 = \a[10][14] ;
    assign _175 = \a[10][15] ;
    assign _176 = \a[11][0] ;
    assign _177 = \a[11][1] ;
    assign _178 = \a[11][2] ;
    assign _179 = \a[11][3] ;
    assign _180 = \a[11][4] ;
    assign _181 = \a[11][5] ;
    assign _182 = \a[11][6] ;
    assign _183 = \a[11][7] ;
    assign _184 = \a[11][8] ;
    assign _185 = \a[11][9] ;
    assign _186 = \a[11][10] ;
    assign _187 = \a[11][11] ;
    assign _188 = \a[11][12] ;
    assign _189 = \a[11][13] ;
    assign _190 = \a[11][14] ;
    assign _191 = \a[11][15] ;
    assign _192 = \a[12][0] ;
    assign _193 = \a[12][1] ;
    assign _194 = \a[12][2] ;
    assign _195 = \a[12][3] ;
    assign _196 = \a[12][4] ;
    assign _197 = \a[12][5] ;
    assign _198 = \a[12][6] ;
    assign _199 = \a[12][7] ;
    assign _200 = \a[12][8] ;
    assign _201 = \a[12][9] ;
    assign _202 = \a[12][10] ;
    assign _203 = \a[12][11] ;
    assign _204 = \a[12][12] ;
    assign _205 = \a[12][13] ;
    assign _206 = \a[12][14] ;
    assign _207 = \a[12][15] ;
    assign _208 = \a[13][0] ;
    assign _209 = \a[13][1] ;
    assign _210 = \a[13][2] ;
    assign _211 = \a[13][3] ;
    assign _212 = \a[13][4] ;
    assign _213 = \a[13][5] ;
    assign _214 = \a[13][6] ;
    assign _215 = \a[13][7] ;
    assign _216 = \a[13][8] ;
    assign _217 = \a[13][9] ;
    assign _218 = \a[13][10] ;
    assign _219 = \a[13][11] ;
    assign _220 = \a[13][12] ;
    assign _221 = \a[13][13] ;
    assign _222 = \a[13][14] ;
    assign _223 = \a[13][15] ;
    assign _224 = \a[14][0] ;
    assign _225 = \a[14][1] ;
    assign _226 = \a[14][2] ;
    assign _227 = \a[14][3] ;
    assign _228 = \a[14][4] ;
    assign _229 = \a[14][5] ;
    assign _230 = \a[14][6] ;
    assign _231 = \a[14][7] ;
    assign _232 = \a[14][8] ;
    assign _233 = \a[14][9] ;
    assign _234 = \a[14][10] ;
    assign _235 = \a[14][11] ;
    assign _236 = \a[14][12] ;
    assign _237 = \a[14][13] ;
    assign _238 = \a[14][14] ;
    assign _239 = \a[14][15] ;
    assign _240 = \a[15][0] ;
    assign _241 = \a[15][1] ;
    assign _242 = \a[15][2] ;
    assign _243 = \a[15][3] ;
    assign _244 = \a[15][4] ;
    assign _245 = \a[15][5] ;
    assign _246 = \a[15][6] ;
    assign _247 = \a[15][7] ;
    assign _248 = \a[15][8] ;
    assign _249 = \a[15][9] ;
    assign _250 = \a[15][10] ;
    assign _251 = \a[15][11] ;
    assign _252 = \a[15][12] ;
    assign _253 = \a[15][13] ;
    assign _254 = \a[15][14] ;
    assign _255 = \a[15][15] ;
    assign \a_sorted[0][0]_ns  = _4319;
    assign \a_sorted[0][1]_ns  = _4320;
    assign \a_sorted[0][2]_ns  = _4321;
    assign \a_sorted[0][3]_ns  = _4322;
    assign \a_sorted[0][4]_ns  = _4323;
    assign \a_sorted[0][5]_ns  = _4324;
    assign \a_sorted[0][6]_ns  = _4325;
    assign \a_sorted[0][7]_ns  = _4326;
    assign \a_sorted[0][8]_ns  = _4327;
    assign \a_sorted[0][9]_ns  = _4328;
    assign \a_sorted[0][10]_ns  = _4329;
    assign \a_sorted[0][11]_ns  = _4330;
    assign \a_sorted[0][12]_ns  = _4331;
    assign \a_sorted[0][13]_ns  = _4332;
    assign \a_sorted[0][14]_ns  = _4333;
    assign \a_sorted[0][15]_ns  = _4334;
    assign \a_sorted[1][0]_ns  = _4335;
    assign \a_sorted[1][1]_ns  = _4336;
    assign \a_sorted[1][2]_ns  = _4337;
    assign \a_sorted[1][3]_ns  = _4338;
    assign \a_sorted[1][4]_ns  = _4339;
    assign \a_sorted[1][5]_ns  = _4340;
    assign \a_sorted[1][6]_ns  = _4341;
    assign \a_sorted[1][7]_ns  = _4342;
    assign \a_sorted[1][8]_ns  = _4343;
    assign \a_sorted[1][9]_ns  = _4344;
    assign \a_sorted[1][10]_ns  = _4345;
    assign \a_sorted[1][11]_ns  = _4346;
    assign \a_sorted[1][12]_ns  = _4347;
    assign \a_sorted[1][13]_ns  = _4348;
    assign \a_sorted[1][14]_ns  = _4349;
    assign \a_sorted[1][15]_ns  = _4350;
    assign \a_sorted[2][0]_ns  = _4384;
    assign \a_sorted[2][1]_ns  = _4385;
    assign \a_sorted[2][2]_ns  = _4386;
    assign \a_sorted[2][3]_ns  = _4387;
    assign \a_sorted[2][4]_ns  = _4388;
    assign \a_sorted[2][5]_ns  = _4389;
    assign \a_sorted[2][6]_ns  = _4390;
    assign \a_sorted[2][7]_ns  = _4391;
    assign \a_sorted[2][8]_ns  = _4392;
    assign \a_sorted[2][9]_ns  = _4393;
    assign \a_sorted[2][10]_ns  = _4394;
    assign \a_sorted[2][11]_ns  = _4395;
    assign \a_sorted[2][12]_ns  = _4396;
    assign \a_sorted[2][13]_ns  = _4397;
    assign \a_sorted[2][14]_ns  = _4398;
    assign \a_sorted[2][15]_ns  = _4399;
    assign \a_sorted[3][0]_ns  = _4400;
    assign \a_sorted[3][1]_ns  = _4401;
    assign \a_sorted[3][2]_ns  = _4402;
    assign \a_sorted[3][3]_ns  = _4403;
    assign \a_sorted[3][4]_ns  = _4404;
    assign \a_sorted[3][5]_ns  = _4405;
    assign \a_sorted[3][6]_ns  = _4406;
    assign \a_sorted[3][7]_ns  = _4407;
    assign \a_sorted[3][8]_ns  = _4408;
    assign \a_sorted[3][9]_ns  = _4409;
    assign \a_sorted[3][10]_ns  = _4410;
    assign \a_sorted[3][11]_ns  = _4411;
    assign \a_sorted[3][12]_ns  = _4412;
    assign \a_sorted[3][13]_ns  = _4413;
    assign \a_sorted[3][14]_ns  = _4414;
    assign \a_sorted[3][15]_ns  = _4415;
    assign \a_sorted[4][0]_ns  = _4579;
    assign \a_sorted[4][1]_ns  = _4580;
    assign \a_sorted[4][2]_ns  = _4581;
    assign \a_sorted[4][3]_ns  = _4582;
    assign \a_sorted[4][4]_ns  = _4583;
    assign \a_sorted[4][5]_ns  = _4584;
    assign \a_sorted[4][6]_ns  = _4585;
    assign \a_sorted[4][7]_ns  = _4586;
    assign \a_sorted[4][8]_ns  = _4587;
    assign \a_sorted[4][9]_ns  = _4588;
    assign \a_sorted[4][10]_ns  = _4589;
    assign \a_sorted[4][11]_ns  = _4590;
    assign \a_sorted[4][12]_ns  = _4591;
    assign \a_sorted[4][13]_ns  = _4592;
    assign \a_sorted[4][14]_ns  = _4593;
    assign \a_sorted[4][15]_ns  = _4594;
    assign \a_sorted[5][0]_ns  = _4595;
    assign \a_sorted[5][1]_ns  = _4596;
    assign \a_sorted[5][2]_ns  = _4597;
    assign \a_sorted[5][3]_ns  = _4598;
    assign \a_sorted[5][4]_ns  = _4599;
    assign \a_sorted[5][5]_ns  = _4600;
    assign \a_sorted[5][6]_ns  = _4601;
    assign \a_sorted[5][7]_ns  = _4602;
    assign \a_sorted[5][8]_ns  = _4603;
    assign \a_sorted[5][9]_ns  = _4604;
    assign \a_sorted[5][10]_ns  = _4605;
    assign \a_sorted[5][11]_ns  = _4606;
    assign \a_sorted[5][12]_ns  = _4607;
    assign \a_sorted[5][13]_ns  = _4608;
    assign \a_sorted[5][14]_ns  = _4609;
    assign \a_sorted[5][15]_ns  = _4610;
    assign \a_sorted[6][0]_ns  = _4644;
    assign \a_sorted[6][1]_ns  = _4645;
    assign \a_sorted[6][2]_ns  = _4646;
    assign \a_sorted[6][3]_ns  = _4647;
    assign \a_sorted[6][4]_ns  = _4648;
    assign \a_sorted[6][5]_ns  = _4649;
    assign \a_sorted[6][6]_ns  = _4650;
    assign \a_sorted[6][7]_ns  = _4651;
    assign \a_sorted[6][8]_ns  = _4652;
    assign \a_sorted[6][9]_ns  = _4653;
    assign \a_sorted[6][10]_ns  = _4654;
    assign \a_sorted[6][11]_ns  = _4655;
    assign \a_sorted[6][12]_ns  = _4656;
    assign \a_sorted[6][13]_ns  = _4657;
    assign \a_sorted[6][14]_ns  = _4658;
    assign \a_sorted[6][15]_ns  = _4659;
    assign \a_sorted[7][0]_ns  = _4660;
    assign \a_sorted[7][1]_ns  = _4661;
    assign \a_sorted[7][2]_ns  = _4662;
    assign \a_sorted[7][3]_ns  = _4663;
    assign \a_sorted[7][4]_ns  = _4664;
    assign \a_sorted[7][5]_ns  = _4665;
    assign \a_sorted[7][6]_ns  = _4666;
    assign \a_sorted[7][7]_ns  = _4667;
    assign \a_sorted[7][8]_ns  = _4668;
    assign \a_sorted[7][9]_ns  = _4669;
    assign \a_sorted[7][10]_ns  = _4670;
    assign \a_sorted[7][11]_ns  = _4671;
    assign \a_sorted[7][12]_ns  = _4672;
    assign \a_sorted[7][13]_ns  = _4673;
    assign \a_sorted[7][14]_ns  = _4674;
    assign \a_sorted[7][15]_ns  = _4675;
    assign \a_sorted[8][0]_ns  = _5099;
    assign \a_sorted[8][1]_ns  = _5100;
    assign \a_sorted[8][2]_ns  = _5101;
    assign \a_sorted[8][3]_ns  = _5102;
    assign \a_sorted[8][4]_ns  = _5103;
    assign \a_sorted[8][5]_ns  = _5104;
    assign \a_sorted[8][6]_ns  = _5105;
    assign \a_sorted[8][7]_ns  = _5106;
    assign \a_sorted[8][8]_ns  = _5107;
    assign \a_sorted[8][9]_ns  = _5108;
    assign \a_sorted[8][10]_ns  = _5109;
    assign \a_sorted[8][11]_ns  = _5110;
    assign \a_sorted[8][12]_ns  = _5111;
    assign \a_sorted[8][13]_ns  = _5112;
    assign \a_sorted[8][14]_ns  = _5113;
    assign \a_sorted[8][15]_ns  = _5114;
    assign \a_sorted[9][0]_ns  = _5115;
    assign \a_sorted[9][1]_ns  = _5116;
    assign \a_sorted[9][2]_ns  = _5117;
    assign \a_sorted[9][3]_ns  = _5118;
    assign \a_sorted[9][4]_ns  = _5119;
    assign \a_sorted[9][5]_ns  = _5120;
    assign \a_sorted[9][6]_ns  = _5121;
    assign \a_sorted[9][7]_ns  = _5122;
    assign \a_sorted[9][8]_ns  = _5123;
    assign \a_sorted[9][9]_ns  = _5124;
    assign \a_sorted[9][10]_ns  = _5125;
    assign \a_sorted[9][11]_ns  = _5126;
    assign \a_sorted[9][12]_ns  = _5127;
    assign \a_sorted[9][13]_ns  = _5128;
    assign \a_sorted[9][14]_ns  = _5129;
    assign \a_sorted[9][15]_ns  = _5130;
    assign \a_sorted[10][0]_ns  = _5164;
    assign \a_sorted[10][1]_ns  = _5165;
    assign \a_sorted[10][2]_ns  = _5166;
    assign \a_sorted[10][3]_ns  = _5167;
    assign \a_sorted[10][4]_ns  = _5168;
    assign \a_sorted[10][5]_ns  = _5169;
    assign \a_sorted[10][6]_ns  = _5170;
    assign \a_sorted[10][7]_ns  = _5171;
    assign \a_sorted[10][8]_ns  = _5172;
    assign \a_sorted[10][9]_ns  = _5173;
    assign \a_sorted[10][10]_ns  = _5174;
    assign \a_sorted[10][11]_ns  = _5175;
    assign \a_sorted[10][12]_ns  = _5176;
    assign \a_sorted[10][13]_ns  = _5177;
    assign \a_sorted[10][14]_ns  = _5178;
    assign \a_sorted[10][15]_ns  = _5179;
    assign \a_sorted[11][0]_ns  = _5180;
    assign \a_sorted[11][1]_ns  = _5181;
    assign \a_sorted[11][2]_ns  = _5182;
    assign \a_sorted[11][3]_ns  = _5183;
    assign \a_sorted[11][4]_ns  = _5184;
    assign \a_sorted[11][5]_ns  = _5185;
    assign \a_sorted[11][6]_ns  = _5186;
    assign \a_sorted[11][7]_ns  = _5187;
    assign \a_sorted[11][8]_ns  = _5188;
    assign \a_sorted[11][9]_ns  = _5189;
    assign \a_sorted[11][10]_ns  = _5190;
    assign \a_sorted[11][11]_ns  = _5191;
    assign \a_sorted[11][12]_ns  = _5192;
    assign \a_sorted[11][13]_ns  = _5193;
    assign \a_sorted[11][14]_ns  = _5194;
    assign \a_sorted[11][15]_ns  = _5195;
    assign \a_sorted[12][0]_ns  = _5359;
    assign \a_sorted[12][1]_ns  = _5360;
    assign \a_sorted[12][2]_ns  = _5361;
    assign \a_sorted[12][3]_ns  = _5362;
    assign \a_sorted[12][4]_ns  = _5363;
    assign \a_sorted[12][5]_ns  = _5364;
    assign \a_sorted[12][6]_ns  = _5365;
    assign \a_sorted[12][7]_ns  = _5366;
    assign \a_sorted[12][8]_ns  = _5367;
    assign \a_sorted[12][9]_ns  = _5368;
    assign \a_sorted[12][10]_ns  = _5369;
    assign \a_sorted[12][11]_ns  = _5370;
    assign \a_sorted[12][12]_ns  = _5371;
    assign \a_sorted[12][13]_ns  = _5372;
    assign \a_sorted[12][14]_ns  = _5373;
    assign \a_sorted[12][15]_ns  = _5374;
    assign \a_sorted[13][0]_ns  = _5375;
    assign \a_sorted[13][1]_ns  = _5376;
    assign \a_sorted[13][2]_ns  = _5377;
    assign \a_sorted[13][3]_ns  = _5378;
    assign \a_sorted[13][4]_ns  = _5379;
    assign \a_sorted[13][5]_ns  = _5380;
    assign \a_sorted[13][6]_ns  = _5381;
    assign \a_sorted[13][7]_ns  = _5382;
    assign \a_sorted[13][8]_ns  = _5383;
    assign \a_sorted[13][9]_ns  = _5384;
    assign \a_sorted[13][10]_ns  = _5385;
    assign \a_sorted[13][11]_ns  = _5386;
    assign \a_sorted[13][12]_ns  = _5387;
    assign \a_sorted[13][13]_ns  = _5388;
    assign \a_sorted[13][14]_ns  = _5389;
    assign \a_sorted[13][15]_ns  = _5390;
    assign \a_sorted[14][0]_ns  = _5424;
    assign \a_sorted[14][1]_ns  = _5425;
    assign \a_sorted[14][2]_ns  = _5426;
    assign \a_sorted[14][3]_ns  = _5427;
    assign \a_sorted[14][4]_ns  = _5428;
    assign \a_sorted[14][5]_ns  = _5429;
    assign \a_sorted[14][6]_ns  = _5430;
    assign \a_sorted[14][7]_ns  = _5431;
    assign \a_sorted[14][8]_ns  = _5432;
    assign \a_sorted[14][9]_ns  = _5433;
    assign \a_sorted[14][10]_ns  = _5434;
    assign \a_sorted[14][11]_ns  = _5435;
    assign \a_sorted[14][12]_ns  = _5436;
    assign \a_sorted[14][13]_ns  = _5437;
    assign \a_sorted[14][14]_ns  = _5438;
    assign \a_sorted[14][15]_ns  = _5439;
    assign \a_sorted[15][0]_ns  = _5440;
    assign \a_sorted[15][1]_ns  = _5441;
    assign \a_sorted[15][2]_ns  = _5442;
    assign \a_sorted[15][3]_ns  = _5443;
    assign \a_sorted[15][4]_ns  = _5444;
    assign \a_sorted[15][5]_ns  = _5445;
    assign \a_sorted[15][6]_ns  = _5446;
    assign \a_sorted[15][7]_ns  = _5447;
    assign \a_sorted[15][8]_ns  = _5448;
    assign \a_sorted[15][9]_ns  = _5449;
    assign \a_sorted[15][10]_ns  = _5450;
    assign \a_sorted[15][11]_ns  = _5451;
    assign \a_sorted[15][12]_ns  = _5452;
    assign \a_sorted[15][13]_ns  = _5453;
    assign \a_sorted[15][14]_ns  = _5454;
    assign \a_sorted[15][15]_ns  = _5455;
    swap u0 (
        .\a[0] (_0),
        .\a[1] (_1),
        .\a[2] (_2),
        .\a[3] (_3),
        .\a[4] (_4),
        .\a[5] (_5),
        .\a[6] (_6),
        .\a[7] (_7),
        .\a[8] (_8),
        .\a[9] (_9),
        .\a[10] (_10),
        .\a[11] (_11),
        .\a[12] (_12),
        .\a[13] (_13),
        .\a[14] (_14),
        .\a[15] (_15),
        .\b[0] (_16),
        .\b[1] (_17),
        .\b[2] (_18),
        .\b[3] (_19),
        .\b[4] (_20),
        .\b[5] (_21),
        .\b[6] (_22),
        .\b[7] (_23),
        .\b[8] (_24),
        .\b[9] (_25),
        .\b[10] (_26),
        .\b[11] (_27),
        .\b[12] (_28),
        .\b[13] (_29),
        .\b[14] (_30),
        .\b[15] (_31),
        .\x[0] (_289),
        .\x[1] (_290),
        .\x[2] (_291),
        .\x[3] (_292),
        .\x[4] (_293),
        .\x[5] (_294),
        .\x[6] (_295),
        .\x[7] (_296),
        .\x[8] (_297),
        .\x[9] (_298),
        .\x[10] (_299),
        .\x[11] (_300),
        .\x[12] (_301),
        .\x[13] (_302),
        .\x[14] (_303),
        .\x[15] (_304),
        .\y[0] (_305),
        .\y[1] (_306),
        .\y[2] (_307),
        .\y[3] (_308),
        .\y[4] (_309),
        .\y[5] (_310),
        .\y[6] (_311),
        .\y[7] (_312),
        .\y[8] (_313),
        .\y[9] (_314),
        .\y[10] (_315),
        .\y[11] (_316),
        .\y[12] (_317),
        .\y[13] (_318),
        .\y[14] (_319),
        .\y[15] (_320)
    );
    swap u1 (
        .\a[0] (_48),
        .\a[1] (_49),
        .\a[2] (_50),
        .\a[3] (_51),
        .\a[4] (_52),
        .\a[5] (_53),
        .\a[6] (_54),
        .\a[7] (_55),
        .\a[8] (_56),
        .\a[9] (_57),
        .\a[10] (_58),
        .\a[11] (_59),
        .\a[12] (_60),
        .\a[13] (_61),
        .\a[14] (_62),
        .\a[15] (_63),
        .\b[0] (_32),
        .\b[1] (_33),
        .\b[2] (_34),
        .\b[3] (_35),
        .\b[4] (_36),
        .\b[5] (_37),
        .\b[6] (_38),
        .\b[7] (_39),
        .\b[8] (_40),
        .\b[9] (_41),
        .\b[10] (_42),
        .\b[11] (_43),
        .\b[12] (_44),
        .\b[13] (_45),
        .\b[14] (_46),
        .\b[15] (_47),
        .\x[0] (_354),
        .\x[1] (_355),
        .\x[2] (_356),
        .\x[3] (_357),
        .\x[4] (_358),
        .\x[5] (_359),
        .\x[6] (_360),
        .\x[7] (_361),
        .\x[8] (_362),
        .\x[9] (_363),
        .\x[10] (_364),
        .\x[11] (_365),
        .\x[12] (_366),
        .\x[13] (_367),
        .\x[14] (_368),
        .\x[15] (_369),
        .\y[0] (_370),
        .\y[1] (_371),
        .\y[2] (_372),
        .\y[3] (_373),
        .\y[4] (_374),
        .\y[5] (_375),
        .\y[6] (_376),
        .\y[7] (_377),
        .\y[8] (_378),
        .\y[9] (_379),
        .\y[10] (_380),
        .\y[11] (_381),
        .\y[12] (_382),
        .\y[13] (_383),
        .\y[14] (_384),
        .\y[15] (_385)
    );
    swap u2 (
        .\a[0] (_289),
        .\a[1] (_290),
        .\a[2] (_291),
        .\a[3] (_292),
        .\a[4] (_293),
        .\a[5] (_294),
        .\a[6] (_295),
        .\a[7] (_296),
        .\a[8] (_297),
        .\a[9] (_298),
        .\a[10] (_299),
        .\a[11] (_300),
        .\a[12] (_301),
        .\a[13] (_302),
        .\a[14] (_303),
        .\a[15] (_304),
        .\b[0] (_370),
        .\b[1] (_371),
        .\b[2] (_372),
        .\b[3] (_373),
        .\b[4] (_374),
        .\b[5] (_375),
        .\b[6] (_376),
        .\b[7] (_377),
        .\b[8] (_378),
        .\b[9] (_379),
        .\b[10] (_380),
        .\b[11] (_381),
        .\b[12] (_382),
        .\b[13] (_383),
        .\b[14] (_384),
        .\b[15] (_385),
        .\x[0] (_419),
        .\x[1] (_420),
        .\x[2] (_421),
        .\x[3] (_422),
        .\x[4] (_423),
        .\x[5] (_424),
        .\x[6] (_425),
        .\x[7] (_426),
        .\x[8] (_427),
        .\x[9] (_428),
        .\x[10] (_429),
        .\x[11] (_430),
        .\x[12] (_431),
        .\x[13] (_432),
        .\x[14] (_433),
        .\x[15] (_434),
        .\y[0] (_435),
        .\y[1] (_436),
        .\y[2] (_437),
        .\y[3] (_438),
        .\y[4] (_439),
        .\y[5] (_440),
        .\y[6] (_441),
        .\y[7] (_442),
        .\y[8] (_443),
        .\y[9] (_444),
        .\y[10] (_445),
        .\y[11] (_446),
        .\y[12] (_447),
        .\y[13] (_448),
        .\y[14] (_449),
        .\y[15] (_450)
    );
    swap u3 (
        .\a[0] (_305),
        .\a[1] (_306),
        .\a[2] (_307),
        .\a[3] (_308),
        .\a[4] (_309),
        .\a[5] (_310),
        .\a[6] (_311),
        .\a[7] (_312),
        .\a[8] (_313),
        .\a[9] (_314),
        .\a[10] (_315),
        .\a[11] (_316),
        .\a[12] (_317),
        .\a[13] (_318),
        .\a[14] (_319),
        .\a[15] (_320),
        .\b[0] (_354),
        .\b[1] (_355),
        .\b[2] (_356),
        .\b[3] (_357),
        .\b[4] (_358),
        .\b[5] (_359),
        .\b[6] (_360),
        .\b[7] (_361),
        .\b[8] (_362),
        .\b[9] (_363),
        .\b[10] (_364),
        .\b[11] (_365),
        .\b[12] (_366),
        .\b[13] (_367),
        .\b[14] (_368),
        .\b[15] (_369),
        .\x[0] (_484),
        .\x[1] (_485),
        .\x[2] (_486),
        .\x[3] (_487),
        .\x[4] (_488),
        .\x[5] (_489),
        .\x[6] (_490),
        .\x[7] (_491),
        .\x[8] (_492),
        .\x[9] (_493),
        .\x[10] (_494),
        .\x[11] (_495),
        .\x[12] (_496),
        .\x[13] (_497),
        .\x[14] (_498),
        .\x[15] (_499),
        .\y[0] (_500),
        .\y[1] (_501),
        .\y[2] (_502),
        .\y[3] (_503),
        .\y[4] (_504),
        .\y[5] (_505),
        .\y[6] (_506),
        .\y[7] (_507),
        .\y[8] (_508),
        .\y[9] (_509),
        .\y[10] (_510),
        .\y[11] (_511),
        .\y[12] (_512),
        .\y[13] (_513),
        .\y[14] (_514),
        .\y[15] (_515)
    );
    swap u4 (
        .\a[0] (_419),
        .\a[1] (_420),
        .\a[2] (_421),
        .\a[3] (_422),
        .\a[4] (_423),
        .\a[5] (_424),
        .\a[6] (_425),
        .\a[7] (_426),
        .\a[8] (_427),
        .\a[9] (_428),
        .\a[10] (_429),
        .\a[11] (_430),
        .\a[12] (_431),
        .\a[13] (_432),
        .\a[14] (_433),
        .\a[15] (_434),
        .\b[0] (_484),
        .\b[1] (_485),
        .\b[2] (_486),
        .\b[3] (_487),
        .\b[4] (_488),
        .\b[5] (_489),
        .\b[6] (_490),
        .\b[7] (_491),
        .\b[8] (_492),
        .\b[9] (_493),
        .\b[10] (_494),
        .\b[11] (_495),
        .\b[12] (_496),
        .\b[13] (_497),
        .\b[14] (_498),
        .\b[15] (_499),
        .\x[0] (_549),
        .\x[1] (_550),
        .\x[2] (_551),
        .\x[3] (_552),
        .\x[4] (_553),
        .\x[5] (_554),
        .\x[6] (_555),
        .\x[7] (_556),
        .\x[8] (_557),
        .\x[9] (_558),
        .\x[10] (_559),
        .\x[11] (_560),
        .\x[12] (_561),
        .\x[13] (_562),
        .\x[14] (_563),
        .\x[15] (_564),
        .\y[0] (_565),
        .\y[1] (_566),
        .\y[2] (_567),
        .\y[3] (_568),
        .\y[4] (_569),
        .\y[5] (_570),
        .\y[6] (_571),
        .\y[7] (_572),
        .\y[8] (_573),
        .\y[9] (_574),
        .\y[10] (_575),
        .\y[11] (_576),
        .\y[12] (_577),
        .\y[13] (_578),
        .\y[14] (_579),
        .\y[15] (_580)
    );
    swap u5 (
        .\a[0] (_435),
        .\a[1] (_436),
        .\a[2] (_437),
        .\a[3] (_438),
        .\a[4] (_439),
        .\a[5] (_440),
        .\a[6] (_441),
        .\a[7] (_442),
        .\a[8] (_443),
        .\a[9] (_444),
        .\a[10] (_445),
        .\a[11] (_446),
        .\a[12] (_447),
        .\a[13] (_448),
        .\a[14] (_449),
        .\a[15] (_450),
        .\b[0] (_500),
        .\b[1] (_501),
        .\b[2] (_502),
        .\b[3] (_503),
        .\b[4] (_504),
        .\b[5] (_505),
        .\b[6] (_506),
        .\b[7] (_507),
        .\b[8] (_508),
        .\b[9] (_509),
        .\b[10] (_510),
        .\b[11] (_511),
        .\b[12] (_512),
        .\b[13] (_513),
        .\b[14] (_514),
        .\b[15] (_515),
        .\x[0] (_614),
        .\x[1] (_615),
        .\x[2] (_616),
        .\x[3] (_617),
        .\x[4] (_618),
        .\x[5] (_619),
        .\x[6] (_620),
        .\x[7] (_621),
        .\x[8] (_622),
        .\x[9] (_623),
        .\x[10] (_624),
        .\x[11] (_625),
        .\x[12] (_626),
        .\x[13] (_627),
        .\x[14] (_628),
        .\x[15] (_629),
        .\y[0] (_630),
        .\y[1] (_631),
        .\y[2] (_632),
        .\y[3] (_633),
        .\y[4] (_634),
        .\y[5] (_635),
        .\y[6] (_636),
        .\y[7] (_637),
        .\y[8] (_638),
        .\y[9] (_639),
        .\y[10] (_640),
        .\y[11] (_641),
        .\y[12] (_642),
        .\y[13] (_643),
        .\y[14] (_644),
        .\y[15] (_645)
    );
    swap u6 (
        .\a[0] (_112),
        .\a[1] (_113),
        .\a[2] (_114),
        .\a[3] (_115),
        .\a[4] (_116),
        .\a[5] (_117),
        .\a[6] (_118),
        .\a[7] (_119),
        .\a[8] (_120),
        .\a[9] (_121),
        .\a[10] (_122),
        .\a[11] (_123),
        .\a[12] (_124),
        .\a[13] (_125),
        .\a[14] (_126),
        .\a[15] (_127),
        .\b[0] (_96),
        .\b[1] (_97),
        .\b[2] (_98),
        .\b[3] (_99),
        .\b[4] (_100),
        .\b[5] (_101),
        .\b[6] (_102),
        .\b[7] (_103),
        .\b[8] (_104),
        .\b[9] (_105),
        .\b[10] (_106),
        .\b[11] (_107),
        .\b[12] (_108),
        .\b[13] (_109),
        .\b[14] (_110),
        .\b[15] (_111),
        .\x[0] (_679),
        .\x[1] (_680),
        .\x[2] (_681),
        .\x[3] (_682),
        .\x[4] (_683),
        .\x[5] (_684),
        .\x[6] (_685),
        .\x[7] (_686),
        .\x[8] (_687),
        .\x[9] (_688),
        .\x[10] (_689),
        .\x[11] (_690),
        .\x[12] (_691),
        .\x[13] (_692),
        .\x[14] (_693),
        .\x[15] (_694),
        .\y[0] (_695),
        .\y[1] (_696),
        .\y[2] (_697),
        .\y[3] (_698),
        .\y[4] (_699),
        .\y[5] (_700),
        .\y[6] (_701),
        .\y[7] (_702),
        .\y[8] (_703),
        .\y[9] (_704),
        .\y[10] (_705),
        .\y[11] (_706),
        .\y[12] (_707),
        .\y[13] (_708),
        .\y[14] (_709),
        .\y[15] (_710)
    );
    swap u7 (
        .\a[0] (_64),
        .\a[1] (_65),
        .\a[2] (_66),
        .\a[3] (_67),
        .\a[4] (_68),
        .\a[5] (_69),
        .\a[6] (_70),
        .\a[7] (_71),
        .\a[8] (_72),
        .\a[9] (_73),
        .\a[10] (_74),
        .\a[11] (_75),
        .\a[12] (_76),
        .\a[13] (_77),
        .\a[14] (_78),
        .\a[15] (_79),
        .\b[0] (_80),
        .\b[1] (_81),
        .\b[2] (_82),
        .\b[3] (_83),
        .\b[4] (_84),
        .\b[5] (_85),
        .\b[6] (_86),
        .\b[7] (_87),
        .\b[8] (_88),
        .\b[9] (_89),
        .\b[10] (_90),
        .\b[11] (_91),
        .\b[12] (_92),
        .\b[13] (_93),
        .\b[14] (_94),
        .\b[15] (_95),
        .\x[0] (_744),
        .\x[1] (_745),
        .\x[2] (_746),
        .\x[3] (_747),
        .\x[4] (_748),
        .\x[5] (_749),
        .\x[6] (_750),
        .\x[7] (_751),
        .\x[8] (_752),
        .\x[9] (_753),
        .\x[10] (_754),
        .\x[11] (_755),
        .\x[12] (_756),
        .\x[13] (_757),
        .\x[14] (_758),
        .\x[15] (_759),
        .\y[0] (_760),
        .\y[1] (_761),
        .\y[2] (_762),
        .\y[3] (_763),
        .\y[4] (_764),
        .\y[5] (_765),
        .\y[6] (_766),
        .\y[7] (_767),
        .\y[8] (_768),
        .\y[9] (_769),
        .\y[10] (_770),
        .\y[11] (_771),
        .\y[12] (_772),
        .\y[13] (_773),
        .\y[14] (_774),
        .\y[15] (_775)
    );
    swap u8 (
        .\a[0] (_679),
        .\a[1] (_680),
        .\a[2] (_681),
        .\a[3] (_682),
        .\a[4] (_683),
        .\a[5] (_684),
        .\a[6] (_685),
        .\a[7] (_686),
        .\a[8] (_687),
        .\a[9] (_688),
        .\a[10] (_689),
        .\a[11] (_690),
        .\a[12] (_691),
        .\a[13] (_692),
        .\a[14] (_693),
        .\a[15] (_694),
        .\b[0] (_760),
        .\b[1] (_761),
        .\b[2] (_762),
        .\b[3] (_763),
        .\b[4] (_764),
        .\b[5] (_765),
        .\b[6] (_766),
        .\b[7] (_767),
        .\b[8] (_768),
        .\b[9] (_769),
        .\b[10] (_770),
        .\b[11] (_771),
        .\b[12] (_772),
        .\b[13] (_773),
        .\b[14] (_774),
        .\b[15] (_775),
        .\x[0] (_809),
        .\x[1] (_810),
        .\x[2] (_811),
        .\x[3] (_812),
        .\x[4] (_813),
        .\x[5] (_814),
        .\x[6] (_815),
        .\x[7] (_816),
        .\x[8] (_817),
        .\x[9] (_818),
        .\x[10] (_819),
        .\x[11] (_820),
        .\x[12] (_821),
        .\x[13] (_822),
        .\x[14] (_823),
        .\x[15] (_824),
        .\y[0] (_825),
        .\y[1] (_826),
        .\y[2] (_827),
        .\y[3] (_828),
        .\y[4] (_829),
        .\y[5] (_830),
        .\y[6] (_831),
        .\y[7] (_832),
        .\y[8] (_833),
        .\y[9] (_834),
        .\y[10] (_835),
        .\y[11] (_836),
        .\y[12] (_837),
        .\y[13] (_838),
        .\y[14] (_839),
        .\y[15] (_840)
    );
    swap u9 (
        .\a[0] (_695),
        .\a[1] (_696),
        .\a[2] (_697),
        .\a[3] (_698),
        .\a[4] (_699),
        .\a[5] (_700),
        .\a[6] (_701),
        .\a[7] (_702),
        .\a[8] (_703),
        .\a[9] (_704),
        .\a[10] (_705),
        .\a[11] (_706),
        .\a[12] (_707),
        .\a[13] (_708),
        .\a[14] (_709),
        .\a[15] (_710),
        .\b[0] (_744),
        .\b[1] (_745),
        .\b[2] (_746),
        .\b[3] (_747),
        .\b[4] (_748),
        .\b[5] (_749),
        .\b[6] (_750),
        .\b[7] (_751),
        .\b[8] (_752),
        .\b[9] (_753),
        .\b[10] (_754),
        .\b[11] (_755),
        .\b[12] (_756),
        .\b[13] (_757),
        .\b[14] (_758),
        .\b[15] (_759),
        .\x[0] (_874),
        .\x[1] (_875),
        .\x[2] (_876),
        .\x[3] (_877),
        .\x[4] (_878),
        .\x[5] (_879),
        .\x[6] (_880),
        .\x[7] (_881),
        .\x[8] (_882),
        .\x[9] (_883),
        .\x[10] (_884),
        .\x[11] (_885),
        .\x[12] (_886),
        .\x[13] (_887),
        .\x[14] (_888),
        .\x[15] (_889),
        .\y[0] (_890),
        .\y[1] (_891),
        .\y[2] (_892),
        .\y[3] (_893),
        .\y[4] (_894),
        .\y[5] (_895),
        .\y[6] (_896),
        .\y[7] (_897),
        .\y[8] (_898),
        .\y[9] (_899),
        .\y[10] (_900),
        .\y[11] (_901),
        .\y[12] (_902),
        .\y[13] (_903),
        .\y[14] (_904),
        .\y[15] (_905)
    );
    swap u10 (
        .\a[0] (_809),
        .\a[1] (_810),
        .\a[2] (_811),
        .\a[3] (_812),
        .\a[4] (_813),
        .\a[5] (_814),
        .\a[6] (_815),
        .\a[7] (_816),
        .\a[8] (_817),
        .\a[9] (_818),
        .\a[10] (_819),
        .\a[11] (_820),
        .\a[12] (_821),
        .\a[13] (_822),
        .\a[14] (_823),
        .\a[15] (_824),
        .\b[0] (_874),
        .\b[1] (_875),
        .\b[2] (_876),
        .\b[3] (_877),
        .\b[4] (_878),
        .\b[5] (_879),
        .\b[6] (_880),
        .\b[7] (_881),
        .\b[8] (_882),
        .\b[9] (_883),
        .\b[10] (_884),
        .\b[11] (_885),
        .\b[12] (_886),
        .\b[13] (_887),
        .\b[14] (_888),
        .\b[15] (_889),
        .\x[0] (_939),
        .\x[1] (_940),
        .\x[2] (_941),
        .\x[3] (_942),
        .\x[4] (_943),
        .\x[5] (_944),
        .\x[6] (_945),
        .\x[7] (_946),
        .\x[8] (_947),
        .\x[9] (_948),
        .\x[10] (_949),
        .\x[11] (_950),
        .\x[12] (_951),
        .\x[13] (_952),
        .\x[14] (_953),
        .\x[15] (_954),
        .\y[0] (_955),
        .\y[1] (_956),
        .\y[2] (_957),
        .\y[3] (_958),
        .\y[4] (_959),
        .\y[5] (_960),
        .\y[6] (_961),
        .\y[7] (_962),
        .\y[8] (_963),
        .\y[9] (_964),
        .\y[10] (_965),
        .\y[11] (_966),
        .\y[12] (_967),
        .\y[13] (_968),
        .\y[14] (_969),
        .\y[15] (_970)
    );
    swap u11 (
        .\a[0] (_825),
        .\a[1] (_826),
        .\a[2] (_827),
        .\a[3] (_828),
        .\a[4] (_829),
        .\a[5] (_830),
        .\a[6] (_831),
        .\a[7] (_832),
        .\a[8] (_833),
        .\a[9] (_834),
        .\a[10] (_835),
        .\a[11] (_836),
        .\a[12] (_837),
        .\a[13] (_838),
        .\a[14] (_839),
        .\a[15] (_840),
        .\b[0] (_890),
        .\b[1] (_891),
        .\b[2] (_892),
        .\b[3] (_893),
        .\b[4] (_894),
        .\b[5] (_895),
        .\b[6] (_896),
        .\b[7] (_897),
        .\b[8] (_898),
        .\b[9] (_899),
        .\b[10] (_900),
        .\b[11] (_901),
        .\b[12] (_902),
        .\b[13] (_903),
        .\b[14] (_904),
        .\b[15] (_905),
        .\x[0] (_1004),
        .\x[1] (_1005),
        .\x[2] (_1006),
        .\x[3] (_1007),
        .\x[4] (_1008),
        .\x[5] (_1009),
        .\x[6] (_1010),
        .\x[7] (_1011),
        .\x[8] (_1012),
        .\x[9] (_1013),
        .\x[10] (_1014),
        .\x[11] (_1015),
        .\x[12] (_1016),
        .\x[13] (_1017),
        .\x[14] (_1018),
        .\x[15] (_1019),
        .\y[0] (_1020),
        .\y[1] (_1021),
        .\y[2] (_1022),
        .\y[3] (_1023),
        .\y[4] (_1024),
        .\y[5] (_1025),
        .\y[6] (_1026),
        .\y[7] (_1027),
        .\y[8] (_1028),
        .\y[9] (_1029),
        .\y[10] (_1030),
        .\y[11] (_1031),
        .\y[12] (_1032),
        .\y[13] (_1033),
        .\y[14] (_1034),
        .\y[15] (_1035)
    );
    swap u12 (
        .\a[0] (_549),
        .\a[1] (_550),
        .\a[2] (_551),
        .\a[3] (_552),
        .\a[4] (_553),
        .\a[5] (_554),
        .\a[6] (_555),
        .\a[7] (_556),
        .\a[8] (_557),
        .\a[9] (_558),
        .\a[10] (_559),
        .\a[11] (_560),
        .\a[12] (_561),
        .\a[13] (_562),
        .\a[14] (_563),
        .\a[15] (_564),
        .\b[0] (_1020),
        .\b[1] (_1021),
        .\b[2] (_1022),
        .\b[3] (_1023),
        .\b[4] (_1024),
        .\b[5] (_1025),
        .\b[6] (_1026),
        .\b[7] (_1027),
        .\b[8] (_1028),
        .\b[9] (_1029),
        .\b[10] (_1030),
        .\b[11] (_1031),
        .\b[12] (_1032),
        .\b[13] (_1033),
        .\b[14] (_1034),
        .\b[15] (_1035),
        .\x[0] (_1069),
        .\x[1] (_1070),
        .\x[2] (_1071),
        .\x[3] (_1072),
        .\x[4] (_1073),
        .\x[5] (_1074),
        .\x[6] (_1075),
        .\x[7] (_1076),
        .\x[8] (_1077),
        .\x[9] (_1078),
        .\x[10] (_1079),
        .\x[11] (_1080),
        .\x[12] (_1081),
        .\x[13] (_1082),
        .\x[14] (_1083),
        .\x[15] (_1084),
        .\y[0] (_1085),
        .\y[1] (_1086),
        .\y[2] (_1087),
        .\y[3] (_1088),
        .\y[4] (_1089),
        .\y[5] (_1090),
        .\y[6] (_1091),
        .\y[7] (_1092),
        .\y[8] (_1093),
        .\y[9] (_1094),
        .\y[10] (_1095),
        .\y[11] (_1096),
        .\y[12] (_1097),
        .\y[13] (_1098),
        .\y[14] (_1099),
        .\y[15] (_1100)
    );
    swap u13 (
        .\a[0] (_565),
        .\a[1] (_566),
        .\a[2] (_567),
        .\a[3] (_568),
        .\a[4] (_569),
        .\a[5] (_570),
        .\a[6] (_571),
        .\a[7] (_572),
        .\a[8] (_573),
        .\a[9] (_574),
        .\a[10] (_575),
        .\a[11] (_576),
        .\a[12] (_577),
        .\a[13] (_578),
        .\a[14] (_579),
        .\a[15] (_580),
        .\b[0] (_1004),
        .\b[1] (_1005),
        .\b[2] (_1006),
        .\b[3] (_1007),
        .\b[4] (_1008),
        .\b[5] (_1009),
        .\b[6] (_1010),
        .\b[7] (_1011),
        .\b[8] (_1012),
        .\b[9] (_1013),
        .\b[10] (_1014),
        .\b[11] (_1015),
        .\b[12] (_1016),
        .\b[13] (_1017),
        .\b[14] (_1018),
        .\b[15] (_1019),
        .\x[0] (_1134),
        .\x[1] (_1135),
        .\x[2] (_1136),
        .\x[3] (_1137),
        .\x[4] (_1138),
        .\x[5] (_1139),
        .\x[6] (_1140),
        .\x[7] (_1141),
        .\x[8] (_1142),
        .\x[9] (_1143),
        .\x[10] (_1144),
        .\x[11] (_1145),
        .\x[12] (_1146),
        .\x[13] (_1147),
        .\x[14] (_1148),
        .\x[15] (_1149),
        .\y[0] (_1150),
        .\y[1] (_1151),
        .\y[2] (_1152),
        .\y[3] (_1153),
        .\y[4] (_1154),
        .\y[5] (_1155),
        .\y[6] (_1156),
        .\y[7] (_1157),
        .\y[8] (_1158),
        .\y[9] (_1159),
        .\y[10] (_1160),
        .\y[11] (_1161),
        .\y[12] (_1162),
        .\y[13] (_1163),
        .\y[14] (_1164),
        .\y[15] (_1165)
    );
    swap u14 (
        .\a[0] (_614),
        .\a[1] (_615),
        .\a[2] (_616),
        .\a[3] (_617),
        .\a[4] (_618),
        .\a[5] (_619),
        .\a[6] (_620),
        .\a[7] (_621),
        .\a[8] (_622),
        .\a[9] (_623),
        .\a[10] (_624),
        .\a[11] (_625),
        .\a[12] (_626),
        .\a[13] (_627),
        .\a[14] (_628),
        .\a[15] (_629),
        .\b[0] (_955),
        .\b[1] (_956),
        .\b[2] (_957),
        .\b[3] (_958),
        .\b[4] (_959),
        .\b[5] (_960),
        .\b[6] (_961),
        .\b[7] (_962),
        .\b[8] (_963),
        .\b[9] (_964),
        .\b[10] (_965),
        .\b[11] (_966),
        .\b[12] (_967),
        .\b[13] (_968),
        .\b[14] (_969),
        .\b[15] (_970),
        .\x[0] (_1199),
        .\x[1] (_1200),
        .\x[2] (_1201),
        .\x[3] (_1202),
        .\x[4] (_1203),
        .\x[5] (_1204),
        .\x[6] (_1205),
        .\x[7] (_1206),
        .\x[8] (_1207),
        .\x[9] (_1208),
        .\x[10] (_1209),
        .\x[11] (_1210),
        .\x[12] (_1211),
        .\x[13] (_1212),
        .\x[14] (_1213),
        .\x[15] (_1214),
        .\y[0] (_1215),
        .\y[1] (_1216),
        .\y[2] (_1217),
        .\y[3] (_1218),
        .\y[4] (_1219),
        .\y[5] (_1220),
        .\y[6] (_1221),
        .\y[7] (_1222),
        .\y[8] (_1223),
        .\y[9] (_1224),
        .\y[10] (_1225),
        .\y[11] (_1226),
        .\y[12] (_1227),
        .\y[13] (_1228),
        .\y[14] (_1229),
        .\y[15] (_1230)
    );
    swap u15 (
        .\a[0] (_630),
        .\a[1] (_631),
        .\a[2] (_632),
        .\a[3] (_633),
        .\a[4] (_634),
        .\a[5] (_635),
        .\a[6] (_636),
        .\a[7] (_637),
        .\a[8] (_638),
        .\a[9] (_639),
        .\a[10] (_640),
        .\a[11] (_641),
        .\a[12] (_642),
        .\a[13] (_643),
        .\a[14] (_644),
        .\a[15] (_645),
        .\b[0] (_939),
        .\b[1] (_940),
        .\b[2] (_941),
        .\b[3] (_942),
        .\b[4] (_943),
        .\b[5] (_944),
        .\b[6] (_945),
        .\b[7] (_946),
        .\b[8] (_947),
        .\b[9] (_948),
        .\b[10] (_949),
        .\b[11] (_950),
        .\b[12] (_951),
        .\b[13] (_952),
        .\b[14] (_953),
        .\b[15] (_954),
        .\x[0] (_1264),
        .\x[1] (_1265),
        .\x[2] (_1266),
        .\x[3] (_1267),
        .\x[4] (_1268),
        .\x[5] (_1269),
        .\x[6] (_1270),
        .\x[7] (_1271),
        .\x[8] (_1272),
        .\x[9] (_1273),
        .\x[10] (_1274),
        .\x[11] (_1275),
        .\x[12] (_1276),
        .\x[13] (_1277),
        .\x[14] (_1278),
        .\x[15] (_1279),
        .\y[0] (_1280),
        .\y[1] (_1281),
        .\y[2] (_1282),
        .\y[3] (_1283),
        .\y[4] (_1284),
        .\y[5] (_1285),
        .\y[6] (_1286),
        .\y[7] (_1287),
        .\y[8] (_1288),
        .\y[9] (_1289),
        .\y[10] (_1290),
        .\y[11] (_1291),
        .\y[12] (_1292),
        .\y[13] (_1293),
        .\y[14] (_1294),
        .\y[15] (_1295)
    );
    swap u16 (
        .\a[0] (_1069),
        .\a[1] (_1070),
        .\a[2] (_1071),
        .\a[3] (_1072),
        .\a[4] (_1073),
        .\a[5] (_1074),
        .\a[6] (_1075),
        .\a[7] (_1076),
        .\a[8] (_1077),
        .\a[9] (_1078),
        .\a[10] (_1079),
        .\a[11] (_1080),
        .\a[12] (_1081),
        .\a[13] (_1082),
        .\a[14] (_1083),
        .\a[15] (_1084),
        .\b[0] (_1199),
        .\b[1] (_1200),
        .\b[2] (_1201),
        .\b[3] (_1202),
        .\b[4] (_1203),
        .\b[5] (_1204),
        .\b[6] (_1205),
        .\b[7] (_1206),
        .\b[8] (_1207),
        .\b[9] (_1208),
        .\b[10] (_1209),
        .\b[11] (_1210),
        .\b[12] (_1211),
        .\b[13] (_1212),
        .\b[14] (_1213),
        .\b[15] (_1214),
        .\x[0] (_1329),
        .\x[1] (_1330),
        .\x[2] (_1331),
        .\x[3] (_1332),
        .\x[4] (_1333),
        .\x[5] (_1334),
        .\x[6] (_1335),
        .\x[7] (_1336),
        .\x[8] (_1337),
        .\x[9] (_1338),
        .\x[10] (_1339),
        .\x[11] (_1340),
        .\x[12] (_1341),
        .\x[13] (_1342),
        .\x[14] (_1343),
        .\x[15] (_1344),
        .\y[0] (_1345),
        .\y[1] (_1346),
        .\y[2] (_1347),
        .\y[3] (_1348),
        .\y[4] (_1349),
        .\y[5] (_1350),
        .\y[6] (_1351),
        .\y[7] (_1352),
        .\y[8] (_1353),
        .\y[9] (_1354),
        .\y[10] (_1355),
        .\y[11] (_1356),
        .\y[12] (_1357),
        .\y[13] (_1358),
        .\y[14] (_1359),
        .\y[15] (_1360)
    );
    swap u17 (
        .\a[0] (_1134),
        .\a[1] (_1135),
        .\a[2] (_1136),
        .\a[3] (_1137),
        .\a[4] (_1138),
        .\a[5] (_1139),
        .\a[6] (_1140),
        .\a[7] (_1141),
        .\a[8] (_1142),
        .\a[9] (_1143),
        .\a[10] (_1144),
        .\a[11] (_1145),
        .\a[12] (_1146),
        .\a[13] (_1147),
        .\a[14] (_1148),
        .\a[15] (_1149),
        .\b[0] (_1264),
        .\b[1] (_1265),
        .\b[2] (_1266),
        .\b[3] (_1267),
        .\b[4] (_1268),
        .\b[5] (_1269),
        .\b[6] (_1270),
        .\b[7] (_1271),
        .\b[8] (_1272),
        .\b[9] (_1273),
        .\b[10] (_1274),
        .\b[11] (_1275),
        .\b[12] (_1276),
        .\b[13] (_1277),
        .\b[14] (_1278),
        .\b[15] (_1279),
        .\x[0] (_1394),
        .\x[1] (_1395),
        .\x[2] (_1396),
        .\x[3] (_1397),
        .\x[4] (_1398),
        .\x[5] (_1399),
        .\x[6] (_1400),
        .\x[7] (_1401),
        .\x[8] (_1402),
        .\x[9] (_1403),
        .\x[10] (_1404),
        .\x[11] (_1405),
        .\x[12] (_1406),
        .\x[13] (_1407),
        .\x[14] (_1408),
        .\x[15] (_1409),
        .\y[0] (_1410),
        .\y[1] (_1411),
        .\y[2] (_1412),
        .\y[3] (_1413),
        .\y[4] (_1414),
        .\y[5] (_1415),
        .\y[6] (_1416),
        .\y[7] (_1417),
        .\y[8] (_1418),
        .\y[9] (_1419),
        .\y[10] (_1420),
        .\y[11] (_1421),
        .\y[12] (_1422),
        .\y[13] (_1423),
        .\y[14] (_1424),
        .\y[15] (_1425)
    );
    swap u18 (
        .\a[0] (_1329),
        .\a[1] (_1330),
        .\a[2] (_1331),
        .\a[3] (_1332),
        .\a[4] (_1333),
        .\a[5] (_1334),
        .\a[6] (_1335),
        .\a[7] (_1336),
        .\a[8] (_1337),
        .\a[9] (_1338),
        .\a[10] (_1339),
        .\a[11] (_1340),
        .\a[12] (_1341),
        .\a[13] (_1342),
        .\a[14] (_1343),
        .\a[15] (_1344),
        .\b[0] (_1394),
        .\b[1] (_1395),
        .\b[2] (_1396),
        .\b[3] (_1397),
        .\b[4] (_1398),
        .\b[5] (_1399),
        .\b[6] (_1400),
        .\b[7] (_1401),
        .\b[8] (_1402),
        .\b[9] (_1403),
        .\b[10] (_1404),
        .\b[11] (_1405),
        .\b[12] (_1406),
        .\b[13] (_1407),
        .\b[14] (_1408),
        .\b[15] (_1409),
        .\x[0] (_1459),
        .\x[1] (_1460),
        .\x[2] (_1461),
        .\x[3] (_1462),
        .\x[4] (_1463),
        .\x[5] (_1464),
        .\x[6] (_1465),
        .\x[7] (_1466),
        .\x[8] (_1467),
        .\x[9] (_1468),
        .\x[10] (_1469),
        .\x[11] (_1470),
        .\x[12] (_1471),
        .\x[13] (_1472),
        .\x[14] (_1473),
        .\x[15] (_1474),
        .\y[0] (_1475),
        .\y[1] (_1476),
        .\y[2] (_1477),
        .\y[3] (_1478),
        .\y[4] (_1479),
        .\y[5] (_1480),
        .\y[6] (_1481),
        .\y[7] (_1482),
        .\y[8] (_1483),
        .\y[9] (_1484),
        .\y[10] (_1485),
        .\y[11] (_1486),
        .\y[12] (_1487),
        .\y[13] (_1488),
        .\y[14] (_1489),
        .\y[15] (_1490)
    );
    swap u19 (
        .\a[0] (_1345),
        .\a[1] (_1346),
        .\a[2] (_1347),
        .\a[3] (_1348),
        .\a[4] (_1349),
        .\a[5] (_1350),
        .\a[6] (_1351),
        .\a[7] (_1352),
        .\a[8] (_1353),
        .\a[9] (_1354),
        .\a[10] (_1355),
        .\a[11] (_1356),
        .\a[12] (_1357),
        .\a[13] (_1358),
        .\a[14] (_1359),
        .\a[15] (_1360),
        .\b[0] (_1410),
        .\b[1] (_1411),
        .\b[2] (_1412),
        .\b[3] (_1413),
        .\b[4] (_1414),
        .\b[5] (_1415),
        .\b[6] (_1416),
        .\b[7] (_1417),
        .\b[8] (_1418),
        .\b[9] (_1419),
        .\b[10] (_1420),
        .\b[11] (_1421),
        .\b[12] (_1422),
        .\b[13] (_1423),
        .\b[14] (_1424),
        .\b[15] (_1425),
        .\x[0] (_1524),
        .\x[1] (_1525),
        .\x[2] (_1526),
        .\x[3] (_1527),
        .\x[4] (_1528),
        .\x[5] (_1529),
        .\x[6] (_1530),
        .\x[7] (_1531),
        .\x[8] (_1532),
        .\x[9] (_1533),
        .\x[10] (_1534),
        .\x[11] (_1535),
        .\x[12] (_1536),
        .\x[13] (_1537),
        .\x[14] (_1538),
        .\x[15] (_1539),
        .\y[0] (_1540),
        .\y[1] (_1541),
        .\y[2] (_1542),
        .\y[3] (_1543),
        .\y[4] (_1544),
        .\y[5] (_1545),
        .\y[6] (_1546),
        .\y[7] (_1547),
        .\y[8] (_1548),
        .\y[9] (_1549),
        .\y[10] (_1550),
        .\y[11] (_1551),
        .\y[12] (_1552),
        .\y[13] (_1553),
        .\y[14] (_1554),
        .\y[15] (_1555)
    );
    swap u20 (
        .\a[0] (_1085),
        .\a[1] (_1086),
        .\a[2] (_1087),
        .\a[3] (_1088),
        .\a[4] (_1089),
        .\a[5] (_1090),
        .\a[6] (_1091),
        .\a[7] (_1092),
        .\a[8] (_1093),
        .\a[9] (_1094),
        .\a[10] (_1095),
        .\a[11] (_1096),
        .\a[12] (_1097),
        .\a[13] (_1098),
        .\a[14] (_1099),
        .\a[15] (_1100),
        .\b[0] (_1215),
        .\b[1] (_1216),
        .\b[2] (_1217),
        .\b[3] (_1218),
        .\b[4] (_1219),
        .\b[5] (_1220),
        .\b[6] (_1221),
        .\b[7] (_1222),
        .\b[8] (_1223),
        .\b[9] (_1224),
        .\b[10] (_1225),
        .\b[11] (_1226),
        .\b[12] (_1227),
        .\b[13] (_1228),
        .\b[14] (_1229),
        .\b[15] (_1230),
        .\x[0] (_1589),
        .\x[1] (_1590),
        .\x[2] (_1591),
        .\x[3] (_1592),
        .\x[4] (_1593),
        .\x[5] (_1594),
        .\x[6] (_1595),
        .\x[7] (_1596),
        .\x[8] (_1597),
        .\x[9] (_1598),
        .\x[10] (_1599),
        .\x[11] (_1600),
        .\x[12] (_1601),
        .\x[13] (_1602),
        .\x[14] (_1603),
        .\x[15] (_1604),
        .\y[0] (_1605),
        .\y[1] (_1606),
        .\y[2] (_1607),
        .\y[3] (_1608),
        .\y[4] (_1609),
        .\y[5] (_1610),
        .\y[6] (_1611),
        .\y[7] (_1612),
        .\y[8] (_1613),
        .\y[9] (_1614),
        .\y[10] (_1615),
        .\y[11] (_1616),
        .\y[12] (_1617),
        .\y[13] (_1618),
        .\y[14] (_1619),
        .\y[15] (_1620)
    );
    swap u21 (
        .\a[0] (_1150),
        .\a[1] (_1151),
        .\a[2] (_1152),
        .\a[3] (_1153),
        .\a[4] (_1154),
        .\a[5] (_1155),
        .\a[6] (_1156),
        .\a[7] (_1157),
        .\a[8] (_1158),
        .\a[9] (_1159),
        .\a[10] (_1160),
        .\a[11] (_1161),
        .\a[12] (_1162),
        .\a[13] (_1163),
        .\a[14] (_1164),
        .\a[15] (_1165),
        .\b[0] (_1280),
        .\b[1] (_1281),
        .\b[2] (_1282),
        .\b[3] (_1283),
        .\b[4] (_1284),
        .\b[5] (_1285),
        .\b[6] (_1286),
        .\b[7] (_1287),
        .\b[8] (_1288),
        .\b[9] (_1289),
        .\b[10] (_1290),
        .\b[11] (_1291),
        .\b[12] (_1292),
        .\b[13] (_1293),
        .\b[14] (_1294),
        .\b[15] (_1295),
        .\x[0] (_1654),
        .\x[1] (_1655),
        .\x[2] (_1656),
        .\x[3] (_1657),
        .\x[4] (_1658),
        .\x[5] (_1659),
        .\x[6] (_1660),
        .\x[7] (_1661),
        .\x[8] (_1662),
        .\x[9] (_1663),
        .\x[10] (_1664),
        .\x[11] (_1665),
        .\x[12] (_1666),
        .\x[13] (_1667),
        .\x[14] (_1668),
        .\x[15] (_1669),
        .\y[0] (_1670),
        .\y[1] (_1671),
        .\y[2] (_1672),
        .\y[3] (_1673),
        .\y[4] (_1674),
        .\y[5] (_1675),
        .\y[6] (_1676),
        .\y[7] (_1677),
        .\y[8] (_1678),
        .\y[9] (_1679),
        .\y[10] (_1680),
        .\y[11] (_1681),
        .\y[12] (_1682),
        .\y[13] (_1683),
        .\y[14] (_1684),
        .\y[15] (_1685)
    );
    swap u22 (
        .\a[0] (_1589),
        .\a[1] (_1590),
        .\a[2] (_1591),
        .\a[3] (_1592),
        .\a[4] (_1593),
        .\a[5] (_1594),
        .\a[6] (_1595),
        .\a[7] (_1596),
        .\a[8] (_1597),
        .\a[9] (_1598),
        .\a[10] (_1599),
        .\a[11] (_1600),
        .\a[12] (_1601),
        .\a[13] (_1602),
        .\a[14] (_1603),
        .\a[15] (_1604),
        .\b[0] (_1654),
        .\b[1] (_1655),
        .\b[2] (_1656),
        .\b[3] (_1657),
        .\b[4] (_1658),
        .\b[5] (_1659),
        .\b[6] (_1660),
        .\b[7] (_1661),
        .\b[8] (_1662),
        .\b[9] (_1663),
        .\b[10] (_1664),
        .\b[11] (_1665),
        .\b[12] (_1666),
        .\b[13] (_1667),
        .\b[14] (_1668),
        .\b[15] (_1669),
        .\x[0] (_1719),
        .\x[1] (_1720),
        .\x[2] (_1721),
        .\x[3] (_1722),
        .\x[4] (_1723),
        .\x[5] (_1724),
        .\x[6] (_1725),
        .\x[7] (_1726),
        .\x[8] (_1727),
        .\x[9] (_1728),
        .\x[10] (_1729),
        .\x[11] (_1730),
        .\x[12] (_1731),
        .\x[13] (_1732),
        .\x[14] (_1733),
        .\x[15] (_1734),
        .\y[0] (_1735),
        .\y[1] (_1736),
        .\y[2] (_1737),
        .\y[3] (_1738),
        .\y[4] (_1739),
        .\y[5] (_1740),
        .\y[6] (_1741),
        .\y[7] (_1742),
        .\y[8] (_1743),
        .\y[9] (_1744),
        .\y[10] (_1745),
        .\y[11] (_1746),
        .\y[12] (_1747),
        .\y[13] (_1748),
        .\y[14] (_1749),
        .\y[15] (_1750)
    );
    swap u23 (
        .\a[0] (_1605),
        .\a[1] (_1606),
        .\a[2] (_1607),
        .\a[3] (_1608),
        .\a[4] (_1609),
        .\a[5] (_1610),
        .\a[6] (_1611),
        .\a[7] (_1612),
        .\a[8] (_1613),
        .\a[9] (_1614),
        .\a[10] (_1615),
        .\a[11] (_1616),
        .\a[12] (_1617),
        .\a[13] (_1618),
        .\a[14] (_1619),
        .\a[15] (_1620),
        .\b[0] (_1670),
        .\b[1] (_1671),
        .\b[2] (_1672),
        .\b[3] (_1673),
        .\b[4] (_1674),
        .\b[5] (_1675),
        .\b[6] (_1676),
        .\b[7] (_1677),
        .\b[8] (_1678),
        .\b[9] (_1679),
        .\b[10] (_1680),
        .\b[11] (_1681),
        .\b[12] (_1682),
        .\b[13] (_1683),
        .\b[14] (_1684),
        .\b[15] (_1685),
        .\x[0] (_1784),
        .\x[1] (_1785),
        .\x[2] (_1786),
        .\x[3] (_1787),
        .\x[4] (_1788),
        .\x[5] (_1789),
        .\x[6] (_1790),
        .\x[7] (_1791),
        .\x[8] (_1792),
        .\x[9] (_1793),
        .\x[10] (_1794),
        .\x[11] (_1795),
        .\x[12] (_1796),
        .\x[13] (_1797),
        .\x[14] (_1798),
        .\x[15] (_1799),
        .\y[0] (_1800),
        .\y[1] (_1801),
        .\y[2] (_1802),
        .\y[3] (_1803),
        .\y[4] (_1804),
        .\y[5] (_1805),
        .\y[6] (_1806),
        .\y[7] (_1807),
        .\y[8] (_1808),
        .\y[9] (_1809),
        .\y[10] (_1810),
        .\y[11] (_1811),
        .\y[12] (_1812),
        .\y[13] (_1813),
        .\y[14] (_1814),
        .\y[15] (_1815)
    );
    swap u24 (
        .\a[0] (_240),
        .\a[1] (_241),
        .\a[2] (_242),
        .\a[3] (_243),
        .\a[4] (_244),
        .\a[5] (_245),
        .\a[6] (_246),
        .\a[7] (_247),
        .\a[8] (_248),
        .\a[9] (_249),
        .\a[10] (_250),
        .\a[11] (_251),
        .\a[12] (_252),
        .\a[13] (_253),
        .\a[14] (_254),
        .\a[15] (_255),
        .\b[0] (_224),
        .\b[1] (_225),
        .\b[2] (_226),
        .\b[3] (_227),
        .\b[4] (_228),
        .\b[5] (_229),
        .\b[6] (_230),
        .\b[7] (_231),
        .\b[8] (_232),
        .\b[9] (_233),
        .\b[10] (_234),
        .\b[11] (_235),
        .\b[12] (_236),
        .\b[13] (_237),
        .\b[14] (_238),
        .\b[15] (_239),
        .\x[0] (_1849),
        .\x[1] (_1850),
        .\x[2] (_1851),
        .\x[3] (_1852),
        .\x[4] (_1853),
        .\x[5] (_1854),
        .\x[6] (_1855),
        .\x[7] (_1856),
        .\x[8] (_1857),
        .\x[9] (_1858),
        .\x[10] (_1859),
        .\x[11] (_1860),
        .\x[12] (_1861),
        .\x[13] (_1862),
        .\x[14] (_1863),
        .\x[15] (_1864),
        .\y[0] (_1865),
        .\y[1] (_1866),
        .\y[2] (_1867),
        .\y[3] (_1868),
        .\y[4] (_1869),
        .\y[5] (_1870),
        .\y[6] (_1871),
        .\y[7] (_1872),
        .\y[8] (_1873),
        .\y[9] (_1874),
        .\y[10] (_1875),
        .\y[11] (_1876),
        .\y[12] (_1877),
        .\y[13] (_1878),
        .\y[14] (_1879),
        .\y[15] (_1880)
    );
    swap u25 (
        .\a[0] (_192),
        .\a[1] (_193),
        .\a[2] (_194),
        .\a[3] (_195),
        .\a[4] (_196),
        .\a[5] (_197),
        .\a[6] (_198),
        .\a[7] (_199),
        .\a[8] (_200),
        .\a[9] (_201),
        .\a[10] (_202),
        .\a[11] (_203),
        .\a[12] (_204),
        .\a[13] (_205),
        .\a[14] (_206),
        .\a[15] (_207),
        .\b[0] (_208),
        .\b[1] (_209),
        .\b[2] (_210),
        .\b[3] (_211),
        .\b[4] (_212),
        .\b[5] (_213),
        .\b[6] (_214),
        .\b[7] (_215),
        .\b[8] (_216),
        .\b[9] (_217),
        .\b[10] (_218),
        .\b[11] (_219),
        .\b[12] (_220),
        .\b[13] (_221),
        .\b[14] (_222),
        .\b[15] (_223),
        .\x[0] (_1914),
        .\x[1] (_1915),
        .\x[2] (_1916),
        .\x[3] (_1917),
        .\x[4] (_1918),
        .\x[5] (_1919),
        .\x[6] (_1920),
        .\x[7] (_1921),
        .\x[8] (_1922),
        .\x[9] (_1923),
        .\x[10] (_1924),
        .\x[11] (_1925),
        .\x[12] (_1926),
        .\x[13] (_1927),
        .\x[14] (_1928),
        .\x[15] (_1929),
        .\y[0] (_1930),
        .\y[1] (_1931),
        .\y[2] (_1932),
        .\y[3] (_1933),
        .\y[4] (_1934),
        .\y[5] (_1935),
        .\y[6] (_1936),
        .\y[7] (_1937),
        .\y[8] (_1938),
        .\y[9] (_1939),
        .\y[10] (_1940),
        .\y[11] (_1941),
        .\y[12] (_1942),
        .\y[13] (_1943),
        .\y[14] (_1944),
        .\y[15] (_1945)
    );
    swap u26 (
        .\a[0] (_1849),
        .\a[1] (_1850),
        .\a[2] (_1851),
        .\a[3] (_1852),
        .\a[4] (_1853),
        .\a[5] (_1854),
        .\a[6] (_1855),
        .\a[7] (_1856),
        .\a[8] (_1857),
        .\a[9] (_1858),
        .\a[10] (_1859),
        .\a[11] (_1860),
        .\a[12] (_1861),
        .\a[13] (_1862),
        .\a[14] (_1863),
        .\a[15] (_1864),
        .\b[0] (_1930),
        .\b[1] (_1931),
        .\b[2] (_1932),
        .\b[3] (_1933),
        .\b[4] (_1934),
        .\b[5] (_1935),
        .\b[6] (_1936),
        .\b[7] (_1937),
        .\b[8] (_1938),
        .\b[9] (_1939),
        .\b[10] (_1940),
        .\b[11] (_1941),
        .\b[12] (_1942),
        .\b[13] (_1943),
        .\b[14] (_1944),
        .\b[15] (_1945),
        .\x[0] (_1979),
        .\x[1] (_1980),
        .\x[2] (_1981),
        .\x[3] (_1982),
        .\x[4] (_1983),
        .\x[5] (_1984),
        .\x[6] (_1985),
        .\x[7] (_1986),
        .\x[8] (_1987),
        .\x[9] (_1988),
        .\x[10] (_1989),
        .\x[11] (_1990),
        .\x[12] (_1991),
        .\x[13] (_1992),
        .\x[14] (_1993),
        .\x[15] (_1994),
        .\y[0] (_1995),
        .\y[1] (_1996),
        .\y[2] (_1997),
        .\y[3] (_1998),
        .\y[4] (_1999),
        .\y[5] (_2000),
        .\y[6] (_2001),
        .\y[7] (_2002),
        .\y[8] (_2003),
        .\y[9] (_2004),
        .\y[10] (_2005),
        .\y[11] (_2006),
        .\y[12] (_2007),
        .\y[13] (_2008),
        .\y[14] (_2009),
        .\y[15] (_2010)
    );
    swap u27 (
        .\a[0] (_1865),
        .\a[1] (_1866),
        .\a[2] (_1867),
        .\a[3] (_1868),
        .\a[4] (_1869),
        .\a[5] (_1870),
        .\a[6] (_1871),
        .\a[7] (_1872),
        .\a[8] (_1873),
        .\a[9] (_1874),
        .\a[10] (_1875),
        .\a[11] (_1876),
        .\a[12] (_1877),
        .\a[13] (_1878),
        .\a[14] (_1879),
        .\a[15] (_1880),
        .\b[0] (_1914),
        .\b[1] (_1915),
        .\b[2] (_1916),
        .\b[3] (_1917),
        .\b[4] (_1918),
        .\b[5] (_1919),
        .\b[6] (_1920),
        .\b[7] (_1921),
        .\b[8] (_1922),
        .\b[9] (_1923),
        .\b[10] (_1924),
        .\b[11] (_1925),
        .\b[12] (_1926),
        .\b[13] (_1927),
        .\b[14] (_1928),
        .\b[15] (_1929),
        .\x[0] (_2044),
        .\x[1] (_2045),
        .\x[2] (_2046),
        .\x[3] (_2047),
        .\x[4] (_2048),
        .\x[5] (_2049),
        .\x[6] (_2050),
        .\x[7] (_2051),
        .\x[8] (_2052),
        .\x[9] (_2053),
        .\x[10] (_2054),
        .\x[11] (_2055),
        .\x[12] (_2056),
        .\x[13] (_2057),
        .\x[14] (_2058),
        .\x[15] (_2059),
        .\y[0] (_2060),
        .\y[1] (_2061),
        .\y[2] (_2062),
        .\y[3] (_2063),
        .\y[4] (_2064),
        .\y[5] (_2065),
        .\y[6] (_2066),
        .\y[7] (_2067),
        .\y[8] (_2068),
        .\y[9] (_2069),
        .\y[10] (_2070),
        .\y[11] (_2071),
        .\y[12] (_2072),
        .\y[13] (_2073),
        .\y[14] (_2074),
        .\y[15] (_2075)
    );
    swap u28 (
        .\a[0] (_1979),
        .\a[1] (_1980),
        .\a[2] (_1981),
        .\a[3] (_1982),
        .\a[4] (_1983),
        .\a[5] (_1984),
        .\a[6] (_1985),
        .\a[7] (_1986),
        .\a[8] (_1987),
        .\a[9] (_1988),
        .\a[10] (_1989),
        .\a[11] (_1990),
        .\a[12] (_1991),
        .\a[13] (_1992),
        .\a[14] (_1993),
        .\a[15] (_1994),
        .\b[0] (_2044),
        .\b[1] (_2045),
        .\b[2] (_2046),
        .\b[3] (_2047),
        .\b[4] (_2048),
        .\b[5] (_2049),
        .\b[6] (_2050),
        .\b[7] (_2051),
        .\b[8] (_2052),
        .\b[9] (_2053),
        .\b[10] (_2054),
        .\b[11] (_2055),
        .\b[12] (_2056),
        .\b[13] (_2057),
        .\b[14] (_2058),
        .\b[15] (_2059),
        .\x[0] (_2109),
        .\x[1] (_2110),
        .\x[2] (_2111),
        .\x[3] (_2112),
        .\x[4] (_2113),
        .\x[5] (_2114),
        .\x[6] (_2115),
        .\x[7] (_2116),
        .\x[8] (_2117),
        .\x[9] (_2118),
        .\x[10] (_2119),
        .\x[11] (_2120),
        .\x[12] (_2121),
        .\x[13] (_2122),
        .\x[14] (_2123),
        .\x[15] (_2124),
        .\y[0] (_2125),
        .\y[1] (_2126),
        .\y[2] (_2127),
        .\y[3] (_2128),
        .\y[4] (_2129),
        .\y[5] (_2130),
        .\y[6] (_2131),
        .\y[7] (_2132),
        .\y[8] (_2133),
        .\y[9] (_2134),
        .\y[10] (_2135),
        .\y[11] (_2136),
        .\y[12] (_2137),
        .\y[13] (_2138),
        .\y[14] (_2139),
        .\y[15] (_2140)
    );
    swap u29 (
        .\a[0] (_1995),
        .\a[1] (_1996),
        .\a[2] (_1997),
        .\a[3] (_1998),
        .\a[4] (_1999),
        .\a[5] (_2000),
        .\a[6] (_2001),
        .\a[7] (_2002),
        .\a[8] (_2003),
        .\a[9] (_2004),
        .\a[10] (_2005),
        .\a[11] (_2006),
        .\a[12] (_2007),
        .\a[13] (_2008),
        .\a[14] (_2009),
        .\a[15] (_2010),
        .\b[0] (_2060),
        .\b[1] (_2061),
        .\b[2] (_2062),
        .\b[3] (_2063),
        .\b[4] (_2064),
        .\b[5] (_2065),
        .\b[6] (_2066),
        .\b[7] (_2067),
        .\b[8] (_2068),
        .\b[9] (_2069),
        .\b[10] (_2070),
        .\b[11] (_2071),
        .\b[12] (_2072),
        .\b[13] (_2073),
        .\b[14] (_2074),
        .\b[15] (_2075),
        .\x[0] (_2174),
        .\x[1] (_2175),
        .\x[2] (_2176),
        .\x[3] (_2177),
        .\x[4] (_2178),
        .\x[5] (_2179),
        .\x[6] (_2180),
        .\x[7] (_2181),
        .\x[8] (_2182),
        .\x[9] (_2183),
        .\x[10] (_2184),
        .\x[11] (_2185),
        .\x[12] (_2186),
        .\x[13] (_2187),
        .\x[14] (_2188),
        .\x[15] (_2189),
        .\y[0] (_2190),
        .\y[1] (_2191),
        .\y[2] (_2192),
        .\y[3] (_2193),
        .\y[4] (_2194),
        .\y[5] (_2195),
        .\y[6] (_2196),
        .\y[7] (_2197),
        .\y[8] (_2198),
        .\y[9] (_2199),
        .\y[10] (_2200),
        .\y[11] (_2201),
        .\y[12] (_2202),
        .\y[13] (_2203),
        .\y[14] (_2204),
        .\y[15] (_2205)
    );
    swap u30 (
        .\a[0] (_128),
        .\a[1] (_129),
        .\a[2] (_130),
        .\a[3] (_131),
        .\a[4] (_132),
        .\a[5] (_133),
        .\a[6] (_134),
        .\a[7] (_135),
        .\a[8] (_136),
        .\a[9] (_137),
        .\a[10] (_138),
        .\a[11] (_139),
        .\a[12] (_140),
        .\a[13] (_141),
        .\a[14] (_142),
        .\a[15] (_143),
        .\b[0] (_144),
        .\b[1] (_145),
        .\b[2] (_146),
        .\b[3] (_147),
        .\b[4] (_148),
        .\b[5] (_149),
        .\b[6] (_150),
        .\b[7] (_151),
        .\b[8] (_152),
        .\b[9] (_153),
        .\b[10] (_154),
        .\b[11] (_155),
        .\b[12] (_156),
        .\b[13] (_157),
        .\b[14] (_158),
        .\b[15] (_159),
        .\x[0] (_2239),
        .\x[1] (_2240),
        .\x[2] (_2241),
        .\x[3] (_2242),
        .\x[4] (_2243),
        .\x[5] (_2244),
        .\x[6] (_2245),
        .\x[7] (_2246),
        .\x[8] (_2247),
        .\x[9] (_2248),
        .\x[10] (_2249),
        .\x[11] (_2250),
        .\x[12] (_2251),
        .\x[13] (_2252),
        .\x[14] (_2253),
        .\x[15] (_2254),
        .\y[0] (_2255),
        .\y[1] (_2256),
        .\y[2] (_2257),
        .\y[3] (_2258),
        .\y[4] (_2259),
        .\y[5] (_2260),
        .\y[6] (_2261),
        .\y[7] (_2262),
        .\y[8] (_2263),
        .\y[9] (_2264),
        .\y[10] (_2265),
        .\y[11] (_2266),
        .\y[12] (_2267),
        .\y[13] (_2268),
        .\y[14] (_2269),
        .\y[15] (_2270)
    );
    swap u31 (
        .\a[0] (_176),
        .\a[1] (_177),
        .\a[2] (_178),
        .\a[3] (_179),
        .\a[4] (_180),
        .\a[5] (_181),
        .\a[6] (_182),
        .\a[7] (_183),
        .\a[8] (_184),
        .\a[9] (_185),
        .\a[10] (_186),
        .\a[11] (_187),
        .\a[12] (_188),
        .\a[13] (_189),
        .\a[14] (_190),
        .\a[15] (_191),
        .\b[0] (_160),
        .\b[1] (_161),
        .\b[2] (_162),
        .\b[3] (_163),
        .\b[4] (_164),
        .\b[5] (_165),
        .\b[6] (_166),
        .\b[7] (_167),
        .\b[8] (_168),
        .\b[9] (_169),
        .\b[10] (_170),
        .\b[11] (_171),
        .\b[12] (_172),
        .\b[13] (_173),
        .\b[14] (_174),
        .\b[15] (_175),
        .\x[0] (_2304),
        .\x[1] (_2305),
        .\x[2] (_2306),
        .\x[3] (_2307),
        .\x[4] (_2308),
        .\x[5] (_2309),
        .\x[6] (_2310),
        .\x[7] (_2311),
        .\x[8] (_2312),
        .\x[9] (_2313),
        .\x[10] (_2314),
        .\x[11] (_2315),
        .\x[12] (_2316),
        .\x[13] (_2317),
        .\x[14] (_2318),
        .\x[15] (_2319),
        .\y[0] (_2320),
        .\y[1] (_2321),
        .\y[2] (_2322),
        .\y[3] (_2323),
        .\y[4] (_2324),
        .\y[5] (_2325),
        .\y[6] (_2326),
        .\y[7] (_2327),
        .\y[8] (_2328),
        .\y[9] (_2329),
        .\y[10] (_2330),
        .\y[11] (_2331),
        .\y[12] (_2332),
        .\y[13] (_2333),
        .\y[14] (_2334),
        .\y[15] (_2335)
    );
    swap u32 (
        .\a[0] (_2239),
        .\a[1] (_2240),
        .\a[2] (_2241),
        .\a[3] (_2242),
        .\a[4] (_2243),
        .\a[5] (_2244),
        .\a[6] (_2245),
        .\a[7] (_2246),
        .\a[8] (_2247),
        .\a[9] (_2248),
        .\a[10] (_2249),
        .\a[11] (_2250),
        .\a[12] (_2251),
        .\a[13] (_2252),
        .\a[14] (_2253),
        .\a[15] (_2254),
        .\b[0] (_2320),
        .\b[1] (_2321),
        .\b[2] (_2322),
        .\b[3] (_2323),
        .\b[4] (_2324),
        .\b[5] (_2325),
        .\b[6] (_2326),
        .\b[7] (_2327),
        .\b[8] (_2328),
        .\b[9] (_2329),
        .\b[10] (_2330),
        .\b[11] (_2331),
        .\b[12] (_2332),
        .\b[13] (_2333),
        .\b[14] (_2334),
        .\b[15] (_2335),
        .\x[0] (_2369),
        .\x[1] (_2370),
        .\x[2] (_2371),
        .\x[3] (_2372),
        .\x[4] (_2373),
        .\x[5] (_2374),
        .\x[6] (_2375),
        .\x[7] (_2376),
        .\x[8] (_2377),
        .\x[9] (_2378),
        .\x[10] (_2379),
        .\x[11] (_2380),
        .\x[12] (_2381),
        .\x[13] (_2382),
        .\x[14] (_2383),
        .\x[15] (_2384),
        .\y[0] (_2385),
        .\y[1] (_2386),
        .\y[2] (_2387),
        .\y[3] (_2388),
        .\y[4] (_2389),
        .\y[5] (_2390),
        .\y[6] (_2391),
        .\y[7] (_2392),
        .\y[8] (_2393),
        .\y[9] (_2394),
        .\y[10] (_2395),
        .\y[11] (_2396),
        .\y[12] (_2397),
        .\y[13] (_2398),
        .\y[14] (_2399),
        .\y[15] (_2400)
    );
    swap u33 (
        .\a[0] (_2255),
        .\a[1] (_2256),
        .\a[2] (_2257),
        .\a[3] (_2258),
        .\a[4] (_2259),
        .\a[5] (_2260),
        .\a[6] (_2261),
        .\a[7] (_2262),
        .\a[8] (_2263),
        .\a[9] (_2264),
        .\a[10] (_2265),
        .\a[11] (_2266),
        .\a[12] (_2267),
        .\a[13] (_2268),
        .\a[14] (_2269),
        .\a[15] (_2270),
        .\b[0] (_2304),
        .\b[1] (_2305),
        .\b[2] (_2306),
        .\b[3] (_2307),
        .\b[4] (_2308),
        .\b[5] (_2309),
        .\b[6] (_2310),
        .\b[7] (_2311),
        .\b[8] (_2312),
        .\b[9] (_2313),
        .\b[10] (_2314),
        .\b[11] (_2315),
        .\b[12] (_2316),
        .\b[13] (_2317),
        .\b[14] (_2318),
        .\b[15] (_2319),
        .\x[0] (_2434),
        .\x[1] (_2435),
        .\x[2] (_2436),
        .\x[3] (_2437),
        .\x[4] (_2438),
        .\x[5] (_2439),
        .\x[6] (_2440),
        .\x[7] (_2441),
        .\x[8] (_2442),
        .\x[9] (_2443),
        .\x[10] (_2444),
        .\x[11] (_2445),
        .\x[12] (_2446),
        .\x[13] (_2447),
        .\x[14] (_2448),
        .\x[15] (_2449),
        .\y[0] (_2450),
        .\y[1] (_2451),
        .\y[2] (_2452),
        .\y[3] (_2453),
        .\y[4] (_2454),
        .\y[5] (_2455),
        .\y[6] (_2456),
        .\y[7] (_2457),
        .\y[8] (_2458),
        .\y[9] (_2459),
        .\y[10] (_2460),
        .\y[11] (_2461),
        .\y[12] (_2462),
        .\y[13] (_2463),
        .\y[14] (_2464),
        .\y[15] (_2465)
    );
    swap u34 (
        .\a[0] (_2369),
        .\a[1] (_2370),
        .\a[2] (_2371),
        .\a[3] (_2372),
        .\a[4] (_2373),
        .\a[5] (_2374),
        .\a[6] (_2375),
        .\a[7] (_2376),
        .\a[8] (_2377),
        .\a[9] (_2378),
        .\a[10] (_2379),
        .\a[11] (_2380),
        .\a[12] (_2381),
        .\a[13] (_2382),
        .\a[14] (_2383),
        .\a[15] (_2384),
        .\b[0] (_2434),
        .\b[1] (_2435),
        .\b[2] (_2436),
        .\b[3] (_2437),
        .\b[4] (_2438),
        .\b[5] (_2439),
        .\b[6] (_2440),
        .\b[7] (_2441),
        .\b[8] (_2442),
        .\b[9] (_2443),
        .\b[10] (_2444),
        .\b[11] (_2445),
        .\b[12] (_2446),
        .\b[13] (_2447),
        .\b[14] (_2448),
        .\b[15] (_2449),
        .\x[0] (_2499),
        .\x[1] (_2500),
        .\x[2] (_2501),
        .\x[3] (_2502),
        .\x[4] (_2503),
        .\x[5] (_2504),
        .\x[6] (_2505),
        .\x[7] (_2506),
        .\x[8] (_2507),
        .\x[9] (_2508),
        .\x[10] (_2509),
        .\x[11] (_2510),
        .\x[12] (_2511),
        .\x[13] (_2512),
        .\x[14] (_2513),
        .\x[15] (_2514),
        .\y[0] (_2515),
        .\y[1] (_2516),
        .\y[2] (_2517),
        .\y[3] (_2518),
        .\y[4] (_2519),
        .\y[5] (_2520),
        .\y[6] (_2521),
        .\y[7] (_2522),
        .\y[8] (_2523),
        .\y[9] (_2524),
        .\y[10] (_2525),
        .\y[11] (_2526),
        .\y[12] (_2527),
        .\y[13] (_2528),
        .\y[14] (_2529),
        .\y[15] (_2530)
    );
    swap u35 (
        .\a[0] (_2385),
        .\a[1] (_2386),
        .\a[2] (_2387),
        .\a[3] (_2388),
        .\a[4] (_2389),
        .\a[5] (_2390),
        .\a[6] (_2391),
        .\a[7] (_2392),
        .\a[8] (_2393),
        .\a[9] (_2394),
        .\a[10] (_2395),
        .\a[11] (_2396),
        .\a[12] (_2397),
        .\a[13] (_2398),
        .\a[14] (_2399),
        .\a[15] (_2400),
        .\b[0] (_2450),
        .\b[1] (_2451),
        .\b[2] (_2452),
        .\b[3] (_2453),
        .\b[4] (_2454),
        .\b[5] (_2455),
        .\b[6] (_2456),
        .\b[7] (_2457),
        .\b[8] (_2458),
        .\b[9] (_2459),
        .\b[10] (_2460),
        .\b[11] (_2461),
        .\b[12] (_2462),
        .\b[13] (_2463),
        .\b[14] (_2464),
        .\b[15] (_2465),
        .\x[0] (_2564),
        .\x[1] (_2565),
        .\x[2] (_2566),
        .\x[3] (_2567),
        .\x[4] (_2568),
        .\x[5] (_2569),
        .\x[6] (_2570),
        .\x[7] (_2571),
        .\x[8] (_2572),
        .\x[9] (_2573),
        .\x[10] (_2574),
        .\x[11] (_2575),
        .\x[12] (_2576),
        .\x[13] (_2577),
        .\x[14] (_2578),
        .\x[15] (_2579),
        .\y[0] (_2580),
        .\y[1] (_2581),
        .\y[2] (_2582),
        .\y[3] (_2583),
        .\y[4] (_2584),
        .\y[5] (_2585),
        .\y[6] (_2586),
        .\y[7] (_2587),
        .\y[8] (_2588),
        .\y[9] (_2589),
        .\y[10] (_2590),
        .\y[11] (_2591),
        .\y[12] (_2592),
        .\y[13] (_2593),
        .\y[14] (_2594),
        .\y[15] (_2595)
    );
    swap u36 (
        .\a[0] (_2109),
        .\a[1] (_2110),
        .\a[2] (_2111),
        .\a[3] (_2112),
        .\a[4] (_2113),
        .\a[5] (_2114),
        .\a[6] (_2115),
        .\a[7] (_2116),
        .\a[8] (_2117),
        .\a[9] (_2118),
        .\a[10] (_2119),
        .\a[11] (_2120),
        .\a[12] (_2121),
        .\a[13] (_2122),
        .\a[14] (_2123),
        .\a[15] (_2124),
        .\b[0] (_2580),
        .\b[1] (_2581),
        .\b[2] (_2582),
        .\b[3] (_2583),
        .\b[4] (_2584),
        .\b[5] (_2585),
        .\b[6] (_2586),
        .\b[7] (_2587),
        .\b[8] (_2588),
        .\b[9] (_2589),
        .\b[10] (_2590),
        .\b[11] (_2591),
        .\b[12] (_2592),
        .\b[13] (_2593),
        .\b[14] (_2594),
        .\b[15] (_2595),
        .\x[0] (_2629),
        .\x[1] (_2630),
        .\x[2] (_2631),
        .\x[3] (_2632),
        .\x[4] (_2633),
        .\x[5] (_2634),
        .\x[6] (_2635),
        .\x[7] (_2636),
        .\x[8] (_2637),
        .\x[9] (_2638),
        .\x[10] (_2639),
        .\x[11] (_2640),
        .\x[12] (_2641),
        .\x[13] (_2642),
        .\x[14] (_2643),
        .\x[15] (_2644),
        .\y[0] (_2645),
        .\y[1] (_2646),
        .\y[2] (_2647),
        .\y[3] (_2648),
        .\y[4] (_2649),
        .\y[5] (_2650),
        .\y[6] (_2651),
        .\y[7] (_2652),
        .\y[8] (_2653),
        .\y[9] (_2654),
        .\y[10] (_2655),
        .\y[11] (_2656),
        .\y[12] (_2657),
        .\y[13] (_2658),
        .\y[14] (_2659),
        .\y[15] (_2660)
    );
    swap u37 (
        .\a[0] (_2125),
        .\a[1] (_2126),
        .\a[2] (_2127),
        .\a[3] (_2128),
        .\a[4] (_2129),
        .\a[5] (_2130),
        .\a[6] (_2131),
        .\a[7] (_2132),
        .\a[8] (_2133),
        .\a[9] (_2134),
        .\a[10] (_2135),
        .\a[11] (_2136),
        .\a[12] (_2137),
        .\a[13] (_2138),
        .\a[14] (_2139),
        .\a[15] (_2140),
        .\b[0] (_2564),
        .\b[1] (_2565),
        .\b[2] (_2566),
        .\b[3] (_2567),
        .\b[4] (_2568),
        .\b[5] (_2569),
        .\b[6] (_2570),
        .\b[7] (_2571),
        .\b[8] (_2572),
        .\b[9] (_2573),
        .\b[10] (_2574),
        .\b[11] (_2575),
        .\b[12] (_2576),
        .\b[13] (_2577),
        .\b[14] (_2578),
        .\b[15] (_2579),
        .\x[0] (_2694),
        .\x[1] (_2695),
        .\x[2] (_2696),
        .\x[3] (_2697),
        .\x[4] (_2698),
        .\x[5] (_2699),
        .\x[6] (_2700),
        .\x[7] (_2701),
        .\x[8] (_2702),
        .\x[9] (_2703),
        .\x[10] (_2704),
        .\x[11] (_2705),
        .\x[12] (_2706),
        .\x[13] (_2707),
        .\x[14] (_2708),
        .\x[15] (_2709),
        .\y[0] (_2710),
        .\y[1] (_2711),
        .\y[2] (_2712),
        .\y[3] (_2713),
        .\y[4] (_2714),
        .\y[5] (_2715),
        .\y[6] (_2716),
        .\y[7] (_2717),
        .\y[8] (_2718),
        .\y[9] (_2719),
        .\y[10] (_2720),
        .\y[11] (_2721),
        .\y[12] (_2722),
        .\y[13] (_2723),
        .\y[14] (_2724),
        .\y[15] (_2725)
    );
    swap u38 (
        .\a[0] (_2174),
        .\a[1] (_2175),
        .\a[2] (_2176),
        .\a[3] (_2177),
        .\a[4] (_2178),
        .\a[5] (_2179),
        .\a[6] (_2180),
        .\a[7] (_2181),
        .\a[8] (_2182),
        .\a[9] (_2183),
        .\a[10] (_2184),
        .\a[11] (_2185),
        .\a[12] (_2186),
        .\a[13] (_2187),
        .\a[14] (_2188),
        .\a[15] (_2189),
        .\b[0] (_2515),
        .\b[1] (_2516),
        .\b[2] (_2517),
        .\b[3] (_2518),
        .\b[4] (_2519),
        .\b[5] (_2520),
        .\b[6] (_2521),
        .\b[7] (_2522),
        .\b[8] (_2523),
        .\b[9] (_2524),
        .\b[10] (_2525),
        .\b[11] (_2526),
        .\b[12] (_2527),
        .\b[13] (_2528),
        .\b[14] (_2529),
        .\b[15] (_2530),
        .\x[0] (_2759),
        .\x[1] (_2760),
        .\x[2] (_2761),
        .\x[3] (_2762),
        .\x[4] (_2763),
        .\x[5] (_2764),
        .\x[6] (_2765),
        .\x[7] (_2766),
        .\x[8] (_2767),
        .\x[9] (_2768),
        .\x[10] (_2769),
        .\x[11] (_2770),
        .\x[12] (_2771),
        .\x[13] (_2772),
        .\x[14] (_2773),
        .\x[15] (_2774),
        .\y[0] (_2775),
        .\y[1] (_2776),
        .\y[2] (_2777),
        .\y[3] (_2778),
        .\y[4] (_2779),
        .\y[5] (_2780),
        .\y[6] (_2781),
        .\y[7] (_2782),
        .\y[8] (_2783),
        .\y[9] (_2784),
        .\y[10] (_2785),
        .\y[11] (_2786),
        .\y[12] (_2787),
        .\y[13] (_2788),
        .\y[14] (_2789),
        .\y[15] (_2790)
    );
    swap u39 (
        .\a[0] (_2190),
        .\a[1] (_2191),
        .\a[2] (_2192),
        .\a[3] (_2193),
        .\a[4] (_2194),
        .\a[5] (_2195),
        .\a[6] (_2196),
        .\a[7] (_2197),
        .\a[8] (_2198),
        .\a[9] (_2199),
        .\a[10] (_2200),
        .\a[11] (_2201),
        .\a[12] (_2202),
        .\a[13] (_2203),
        .\a[14] (_2204),
        .\a[15] (_2205),
        .\b[0] (_2499),
        .\b[1] (_2500),
        .\b[2] (_2501),
        .\b[3] (_2502),
        .\b[4] (_2503),
        .\b[5] (_2504),
        .\b[6] (_2505),
        .\b[7] (_2506),
        .\b[8] (_2507),
        .\b[9] (_2508),
        .\b[10] (_2509),
        .\b[11] (_2510),
        .\b[12] (_2511),
        .\b[13] (_2512),
        .\b[14] (_2513),
        .\b[15] (_2514),
        .\x[0] (_2824),
        .\x[1] (_2825),
        .\x[2] (_2826),
        .\x[3] (_2827),
        .\x[4] (_2828),
        .\x[5] (_2829),
        .\x[6] (_2830),
        .\x[7] (_2831),
        .\x[8] (_2832),
        .\x[9] (_2833),
        .\x[10] (_2834),
        .\x[11] (_2835),
        .\x[12] (_2836),
        .\x[13] (_2837),
        .\x[14] (_2838),
        .\x[15] (_2839),
        .\y[0] (_2840),
        .\y[1] (_2841),
        .\y[2] (_2842),
        .\y[3] (_2843),
        .\y[4] (_2844),
        .\y[5] (_2845),
        .\y[6] (_2846),
        .\y[7] (_2847),
        .\y[8] (_2848),
        .\y[9] (_2849),
        .\y[10] (_2850),
        .\y[11] (_2851),
        .\y[12] (_2852),
        .\y[13] (_2853),
        .\y[14] (_2854),
        .\y[15] (_2855)
    );
    swap u40 (
        .\a[0] (_2629),
        .\a[1] (_2630),
        .\a[2] (_2631),
        .\a[3] (_2632),
        .\a[4] (_2633),
        .\a[5] (_2634),
        .\a[6] (_2635),
        .\a[7] (_2636),
        .\a[8] (_2637),
        .\a[9] (_2638),
        .\a[10] (_2639),
        .\a[11] (_2640),
        .\a[12] (_2641),
        .\a[13] (_2642),
        .\a[14] (_2643),
        .\a[15] (_2644),
        .\b[0] (_2759),
        .\b[1] (_2760),
        .\b[2] (_2761),
        .\b[3] (_2762),
        .\b[4] (_2763),
        .\b[5] (_2764),
        .\b[6] (_2765),
        .\b[7] (_2766),
        .\b[8] (_2767),
        .\b[9] (_2768),
        .\b[10] (_2769),
        .\b[11] (_2770),
        .\b[12] (_2771),
        .\b[13] (_2772),
        .\b[14] (_2773),
        .\b[15] (_2774),
        .\x[0] (_2889),
        .\x[1] (_2890),
        .\x[2] (_2891),
        .\x[3] (_2892),
        .\x[4] (_2893),
        .\x[5] (_2894),
        .\x[6] (_2895),
        .\x[7] (_2896),
        .\x[8] (_2897),
        .\x[9] (_2898),
        .\x[10] (_2899),
        .\x[11] (_2900),
        .\x[12] (_2901),
        .\x[13] (_2902),
        .\x[14] (_2903),
        .\x[15] (_2904),
        .\y[0] (_2905),
        .\y[1] (_2906),
        .\y[2] (_2907),
        .\y[3] (_2908),
        .\y[4] (_2909),
        .\y[5] (_2910),
        .\y[6] (_2911),
        .\y[7] (_2912),
        .\y[8] (_2913),
        .\y[9] (_2914),
        .\y[10] (_2915),
        .\y[11] (_2916),
        .\y[12] (_2917),
        .\y[13] (_2918),
        .\y[14] (_2919),
        .\y[15] (_2920)
    );
    swap u41 (
        .\a[0] (_2694),
        .\a[1] (_2695),
        .\a[2] (_2696),
        .\a[3] (_2697),
        .\a[4] (_2698),
        .\a[5] (_2699),
        .\a[6] (_2700),
        .\a[7] (_2701),
        .\a[8] (_2702),
        .\a[9] (_2703),
        .\a[10] (_2704),
        .\a[11] (_2705),
        .\a[12] (_2706),
        .\a[13] (_2707),
        .\a[14] (_2708),
        .\a[15] (_2709),
        .\b[0] (_2824),
        .\b[1] (_2825),
        .\b[2] (_2826),
        .\b[3] (_2827),
        .\b[4] (_2828),
        .\b[5] (_2829),
        .\b[6] (_2830),
        .\b[7] (_2831),
        .\b[8] (_2832),
        .\b[9] (_2833),
        .\b[10] (_2834),
        .\b[11] (_2835),
        .\b[12] (_2836),
        .\b[13] (_2837),
        .\b[14] (_2838),
        .\b[15] (_2839),
        .\x[0] (_2954),
        .\x[1] (_2955),
        .\x[2] (_2956),
        .\x[3] (_2957),
        .\x[4] (_2958),
        .\x[5] (_2959),
        .\x[6] (_2960),
        .\x[7] (_2961),
        .\x[8] (_2962),
        .\x[9] (_2963),
        .\x[10] (_2964),
        .\x[11] (_2965),
        .\x[12] (_2966),
        .\x[13] (_2967),
        .\x[14] (_2968),
        .\x[15] (_2969),
        .\y[0] (_2970),
        .\y[1] (_2971),
        .\y[2] (_2972),
        .\y[3] (_2973),
        .\y[4] (_2974),
        .\y[5] (_2975),
        .\y[6] (_2976),
        .\y[7] (_2977),
        .\y[8] (_2978),
        .\y[9] (_2979),
        .\y[10] (_2980),
        .\y[11] (_2981),
        .\y[12] (_2982),
        .\y[13] (_2983),
        .\y[14] (_2984),
        .\y[15] (_2985)
    );
    swap u42 (
        .\a[0] (_2889),
        .\a[1] (_2890),
        .\a[2] (_2891),
        .\a[3] (_2892),
        .\a[4] (_2893),
        .\a[5] (_2894),
        .\a[6] (_2895),
        .\a[7] (_2896),
        .\a[8] (_2897),
        .\a[9] (_2898),
        .\a[10] (_2899),
        .\a[11] (_2900),
        .\a[12] (_2901),
        .\a[13] (_2902),
        .\a[14] (_2903),
        .\a[15] (_2904),
        .\b[0] (_2954),
        .\b[1] (_2955),
        .\b[2] (_2956),
        .\b[3] (_2957),
        .\b[4] (_2958),
        .\b[5] (_2959),
        .\b[6] (_2960),
        .\b[7] (_2961),
        .\b[8] (_2962),
        .\b[9] (_2963),
        .\b[10] (_2964),
        .\b[11] (_2965),
        .\b[12] (_2966),
        .\b[13] (_2967),
        .\b[14] (_2968),
        .\b[15] (_2969),
        .\x[0] (_3019),
        .\x[1] (_3020),
        .\x[2] (_3021),
        .\x[3] (_3022),
        .\x[4] (_3023),
        .\x[5] (_3024),
        .\x[6] (_3025),
        .\x[7] (_3026),
        .\x[8] (_3027),
        .\x[9] (_3028),
        .\x[10] (_3029),
        .\x[11] (_3030),
        .\x[12] (_3031),
        .\x[13] (_3032),
        .\x[14] (_3033),
        .\x[15] (_3034),
        .\y[0] (_3035),
        .\y[1] (_3036),
        .\y[2] (_3037),
        .\y[3] (_3038),
        .\y[4] (_3039),
        .\y[5] (_3040),
        .\y[6] (_3041),
        .\y[7] (_3042),
        .\y[8] (_3043),
        .\y[9] (_3044),
        .\y[10] (_3045),
        .\y[11] (_3046),
        .\y[12] (_3047),
        .\y[13] (_3048),
        .\y[14] (_3049),
        .\y[15] (_3050)
    );
    swap u43 (
        .\a[0] (_2905),
        .\a[1] (_2906),
        .\a[2] (_2907),
        .\a[3] (_2908),
        .\a[4] (_2909),
        .\a[5] (_2910),
        .\a[6] (_2911),
        .\a[7] (_2912),
        .\a[8] (_2913),
        .\a[9] (_2914),
        .\a[10] (_2915),
        .\a[11] (_2916),
        .\a[12] (_2917),
        .\a[13] (_2918),
        .\a[14] (_2919),
        .\a[15] (_2920),
        .\b[0] (_2970),
        .\b[1] (_2971),
        .\b[2] (_2972),
        .\b[3] (_2973),
        .\b[4] (_2974),
        .\b[5] (_2975),
        .\b[6] (_2976),
        .\b[7] (_2977),
        .\b[8] (_2978),
        .\b[9] (_2979),
        .\b[10] (_2980),
        .\b[11] (_2981),
        .\b[12] (_2982),
        .\b[13] (_2983),
        .\b[14] (_2984),
        .\b[15] (_2985),
        .\x[0] (_3084),
        .\x[1] (_3085),
        .\x[2] (_3086),
        .\x[3] (_3087),
        .\x[4] (_3088),
        .\x[5] (_3089),
        .\x[6] (_3090),
        .\x[7] (_3091),
        .\x[8] (_3092),
        .\x[9] (_3093),
        .\x[10] (_3094),
        .\x[11] (_3095),
        .\x[12] (_3096),
        .\x[13] (_3097),
        .\x[14] (_3098),
        .\x[15] (_3099),
        .\y[0] (_3100),
        .\y[1] (_3101),
        .\y[2] (_3102),
        .\y[3] (_3103),
        .\y[4] (_3104),
        .\y[5] (_3105),
        .\y[6] (_3106),
        .\y[7] (_3107),
        .\y[8] (_3108),
        .\y[9] (_3109),
        .\y[10] (_3110),
        .\y[11] (_3111),
        .\y[12] (_3112),
        .\y[13] (_3113),
        .\y[14] (_3114),
        .\y[15] (_3115)
    );
    swap u44 (
        .\a[0] (_2645),
        .\a[1] (_2646),
        .\a[2] (_2647),
        .\a[3] (_2648),
        .\a[4] (_2649),
        .\a[5] (_2650),
        .\a[6] (_2651),
        .\a[7] (_2652),
        .\a[8] (_2653),
        .\a[9] (_2654),
        .\a[10] (_2655),
        .\a[11] (_2656),
        .\a[12] (_2657),
        .\a[13] (_2658),
        .\a[14] (_2659),
        .\a[15] (_2660),
        .\b[0] (_2775),
        .\b[1] (_2776),
        .\b[2] (_2777),
        .\b[3] (_2778),
        .\b[4] (_2779),
        .\b[5] (_2780),
        .\b[6] (_2781),
        .\b[7] (_2782),
        .\b[8] (_2783),
        .\b[9] (_2784),
        .\b[10] (_2785),
        .\b[11] (_2786),
        .\b[12] (_2787),
        .\b[13] (_2788),
        .\b[14] (_2789),
        .\b[15] (_2790),
        .\x[0] (_3149),
        .\x[1] (_3150),
        .\x[2] (_3151),
        .\x[3] (_3152),
        .\x[4] (_3153),
        .\x[5] (_3154),
        .\x[6] (_3155),
        .\x[7] (_3156),
        .\x[8] (_3157),
        .\x[9] (_3158),
        .\x[10] (_3159),
        .\x[11] (_3160),
        .\x[12] (_3161),
        .\x[13] (_3162),
        .\x[14] (_3163),
        .\x[15] (_3164),
        .\y[0] (_3165),
        .\y[1] (_3166),
        .\y[2] (_3167),
        .\y[3] (_3168),
        .\y[4] (_3169),
        .\y[5] (_3170),
        .\y[6] (_3171),
        .\y[7] (_3172),
        .\y[8] (_3173),
        .\y[9] (_3174),
        .\y[10] (_3175),
        .\y[11] (_3176),
        .\y[12] (_3177),
        .\y[13] (_3178),
        .\y[14] (_3179),
        .\y[15] (_3180)
    );
    swap u45 (
        .\a[0] (_2710),
        .\a[1] (_2711),
        .\a[2] (_2712),
        .\a[3] (_2713),
        .\a[4] (_2714),
        .\a[5] (_2715),
        .\a[6] (_2716),
        .\a[7] (_2717),
        .\a[8] (_2718),
        .\a[9] (_2719),
        .\a[10] (_2720),
        .\a[11] (_2721),
        .\a[12] (_2722),
        .\a[13] (_2723),
        .\a[14] (_2724),
        .\a[15] (_2725),
        .\b[0] (_2840),
        .\b[1] (_2841),
        .\b[2] (_2842),
        .\b[3] (_2843),
        .\b[4] (_2844),
        .\b[5] (_2845),
        .\b[6] (_2846),
        .\b[7] (_2847),
        .\b[8] (_2848),
        .\b[9] (_2849),
        .\b[10] (_2850),
        .\b[11] (_2851),
        .\b[12] (_2852),
        .\b[13] (_2853),
        .\b[14] (_2854),
        .\b[15] (_2855),
        .\x[0] (_3214),
        .\x[1] (_3215),
        .\x[2] (_3216),
        .\x[3] (_3217),
        .\x[4] (_3218),
        .\x[5] (_3219),
        .\x[6] (_3220),
        .\x[7] (_3221),
        .\x[8] (_3222),
        .\x[9] (_3223),
        .\x[10] (_3224),
        .\x[11] (_3225),
        .\x[12] (_3226),
        .\x[13] (_3227),
        .\x[14] (_3228),
        .\x[15] (_3229),
        .\y[0] (_3230),
        .\y[1] (_3231),
        .\y[2] (_3232),
        .\y[3] (_3233),
        .\y[4] (_3234),
        .\y[5] (_3235),
        .\y[6] (_3236),
        .\y[7] (_3237),
        .\y[8] (_3238),
        .\y[9] (_3239),
        .\y[10] (_3240),
        .\y[11] (_3241),
        .\y[12] (_3242),
        .\y[13] (_3243),
        .\y[14] (_3244),
        .\y[15] (_3245)
    );
    swap u46 (
        .\a[0] (_3149),
        .\a[1] (_3150),
        .\a[2] (_3151),
        .\a[3] (_3152),
        .\a[4] (_3153),
        .\a[5] (_3154),
        .\a[6] (_3155),
        .\a[7] (_3156),
        .\a[8] (_3157),
        .\a[9] (_3158),
        .\a[10] (_3159),
        .\a[11] (_3160),
        .\a[12] (_3161),
        .\a[13] (_3162),
        .\a[14] (_3163),
        .\a[15] (_3164),
        .\b[0] (_3214),
        .\b[1] (_3215),
        .\b[2] (_3216),
        .\b[3] (_3217),
        .\b[4] (_3218),
        .\b[5] (_3219),
        .\b[6] (_3220),
        .\b[7] (_3221),
        .\b[8] (_3222),
        .\b[9] (_3223),
        .\b[10] (_3224),
        .\b[11] (_3225),
        .\b[12] (_3226),
        .\b[13] (_3227),
        .\b[14] (_3228),
        .\b[15] (_3229),
        .\x[0] (_3279),
        .\x[1] (_3280),
        .\x[2] (_3281),
        .\x[3] (_3282),
        .\x[4] (_3283),
        .\x[5] (_3284),
        .\x[6] (_3285),
        .\x[7] (_3286),
        .\x[8] (_3287),
        .\x[9] (_3288),
        .\x[10] (_3289),
        .\x[11] (_3290),
        .\x[12] (_3291),
        .\x[13] (_3292),
        .\x[14] (_3293),
        .\x[15] (_3294),
        .\y[0] (_3295),
        .\y[1] (_3296),
        .\y[2] (_3297),
        .\y[3] (_3298),
        .\y[4] (_3299),
        .\y[5] (_3300),
        .\y[6] (_3301),
        .\y[7] (_3302),
        .\y[8] (_3303),
        .\y[9] (_3304),
        .\y[10] (_3305),
        .\y[11] (_3306),
        .\y[12] (_3307),
        .\y[13] (_3308),
        .\y[14] (_3309),
        .\y[15] (_3310)
    );
    swap u47 (
        .\a[0] (_3165),
        .\a[1] (_3166),
        .\a[2] (_3167),
        .\a[3] (_3168),
        .\a[4] (_3169),
        .\a[5] (_3170),
        .\a[6] (_3171),
        .\a[7] (_3172),
        .\a[8] (_3173),
        .\a[9] (_3174),
        .\a[10] (_3175),
        .\a[11] (_3176),
        .\a[12] (_3177),
        .\a[13] (_3178),
        .\a[14] (_3179),
        .\a[15] (_3180),
        .\b[0] (_3230),
        .\b[1] (_3231),
        .\b[2] (_3232),
        .\b[3] (_3233),
        .\b[4] (_3234),
        .\b[5] (_3235),
        .\b[6] (_3236),
        .\b[7] (_3237),
        .\b[8] (_3238),
        .\b[9] (_3239),
        .\b[10] (_3240),
        .\b[11] (_3241),
        .\b[12] (_3242),
        .\b[13] (_3243),
        .\b[14] (_3244),
        .\b[15] (_3245),
        .\x[0] (_3344),
        .\x[1] (_3345),
        .\x[2] (_3346),
        .\x[3] (_3347),
        .\x[4] (_3348),
        .\x[5] (_3349),
        .\x[6] (_3350),
        .\x[7] (_3351),
        .\x[8] (_3352),
        .\x[9] (_3353),
        .\x[10] (_3354),
        .\x[11] (_3355),
        .\x[12] (_3356),
        .\x[13] (_3357),
        .\x[14] (_3358),
        .\x[15] (_3359),
        .\y[0] (_3360),
        .\y[1] (_3361),
        .\y[2] (_3362),
        .\y[3] (_3363),
        .\y[4] (_3364),
        .\y[5] (_3365),
        .\y[6] (_3366),
        .\y[7] (_3367),
        .\y[8] (_3368),
        .\y[9] (_3369),
        .\y[10] (_3370),
        .\y[11] (_3371),
        .\y[12] (_3372),
        .\y[13] (_3373),
        .\y[14] (_3374),
        .\y[15] (_3375)
    );
    swap u48 (
        .\a[0] (_1459),
        .\a[1] (_1460),
        .\a[2] (_1461),
        .\a[3] (_1462),
        .\a[4] (_1463),
        .\a[5] (_1464),
        .\a[6] (_1465),
        .\a[7] (_1466),
        .\a[8] (_1467),
        .\a[9] (_1468),
        .\a[10] (_1469),
        .\a[11] (_1470),
        .\a[12] (_1471),
        .\a[13] (_1472),
        .\a[14] (_1473),
        .\a[15] (_1474),
        .\b[0] (_3360),
        .\b[1] (_3361),
        .\b[2] (_3362),
        .\b[3] (_3363),
        .\b[4] (_3364),
        .\b[5] (_3365),
        .\b[6] (_3366),
        .\b[7] (_3367),
        .\b[8] (_3368),
        .\b[9] (_3369),
        .\b[10] (_3370),
        .\b[11] (_3371),
        .\b[12] (_3372),
        .\b[13] (_3373),
        .\b[14] (_3374),
        .\b[15] (_3375),
        .\x[0] (_3409),
        .\x[1] (_3410),
        .\x[2] (_3411),
        .\x[3] (_3412),
        .\x[4] (_3413),
        .\x[5] (_3414),
        .\x[6] (_3415),
        .\x[7] (_3416),
        .\x[8] (_3417),
        .\x[9] (_3418),
        .\x[10] (_3419),
        .\x[11] (_3420),
        .\x[12] (_3421),
        .\x[13] (_3422),
        .\x[14] (_3423),
        .\x[15] (_3424),
        .\y[0] (_3425),
        .\y[1] (_3426),
        .\y[2] (_3427),
        .\y[3] (_3428),
        .\y[4] (_3429),
        .\y[5] (_3430),
        .\y[6] (_3431),
        .\y[7] (_3432),
        .\y[8] (_3433),
        .\y[9] (_3434),
        .\y[10] (_3435),
        .\y[11] (_3436),
        .\y[12] (_3437),
        .\y[13] (_3438),
        .\y[14] (_3439),
        .\y[15] (_3440)
    );
    swap u49 (
        .\a[0] (_1475),
        .\a[1] (_1476),
        .\a[2] (_1477),
        .\a[3] (_1478),
        .\a[4] (_1479),
        .\a[5] (_1480),
        .\a[6] (_1481),
        .\a[7] (_1482),
        .\a[8] (_1483),
        .\a[9] (_1484),
        .\a[10] (_1485),
        .\a[11] (_1486),
        .\a[12] (_1487),
        .\a[13] (_1488),
        .\a[14] (_1489),
        .\a[15] (_1490),
        .\b[0] (_3344),
        .\b[1] (_3345),
        .\b[2] (_3346),
        .\b[3] (_3347),
        .\b[4] (_3348),
        .\b[5] (_3349),
        .\b[6] (_3350),
        .\b[7] (_3351),
        .\b[8] (_3352),
        .\b[9] (_3353),
        .\b[10] (_3354),
        .\b[11] (_3355),
        .\b[12] (_3356),
        .\b[13] (_3357),
        .\b[14] (_3358),
        .\b[15] (_3359),
        .\x[0] (_3474),
        .\x[1] (_3475),
        .\x[2] (_3476),
        .\x[3] (_3477),
        .\x[4] (_3478),
        .\x[5] (_3479),
        .\x[6] (_3480),
        .\x[7] (_3481),
        .\x[8] (_3482),
        .\x[9] (_3483),
        .\x[10] (_3484),
        .\x[11] (_3485),
        .\x[12] (_3486),
        .\x[13] (_3487),
        .\x[14] (_3488),
        .\x[15] (_3489),
        .\y[0] (_3490),
        .\y[1] (_3491),
        .\y[2] (_3492),
        .\y[3] (_3493),
        .\y[4] (_3494),
        .\y[5] (_3495),
        .\y[6] (_3496),
        .\y[7] (_3497),
        .\y[8] (_3498),
        .\y[9] (_3499),
        .\y[10] (_3500),
        .\y[11] (_3501),
        .\y[12] (_3502),
        .\y[13] (_3503),
        .\y[14] (_3504),
        .\y[15] (_3505)
    );
    swap u50 (
        .\a[0] (_1524),
        .\a[1] (_1525),
        .\a[2] (_1526),
        .\a[3] (_1527),
        .\a[4] (_1528),
        .\a[5] (_1529),
        .\a[6] (_1530),
        .\a[7] (_1531),
        .\a[8] (_1532),
        .\a[9] (_1533),
        .\a[10] (_1534),
        .\a[11] (_1535),
        .\a[12] (_1536),
        .\a[13] (_1537),
        .\a[14] (_1538),
        .\a[15] (_1539),
        .\b[0] (_3295),
        .\b[1] (_3296),
        .\b[2] (_3297),
        .\b[3] (_3298),
        .\b[4] (_3299),
        .\b[5] (_3300),
        .\b[6] (_3301),
        .\b[7] (_3302),
        .\b[8] (_3303),
        .\b[9] (_3304),
        .\b[10] (_3305),
        .\b[11] (_3306),
        .\b[12] (_3307),
        .\b[13] (_3308),
        .\b[14] (_3309),
        .\b[15] (_3310),
        .\x[0] (_3539),
        .\x[1] (_3540),
        .\x[2] (_3541),
        .\x[3] (_3542),
        .\x[4] (_3543),
        .\x[5] (_3544),
        .\x[6] (_3545),
        .\x[7] (_3546),
        .\x[8] (_3547),
        .\x[9] (_3548),
        .\x[10] (_3549),
        .\x[11] (_3550),
        .\x[12] (_3551),
        .\x[13] (_3552),
        .\x[14] (_3553),
        .\x[15] (_3554),
        .\y[0] (_3555),
        .\y[1] (_3556),
        .\y[2] (_3557),
        .\y[3] (_3558),
        .\y[4] (_3559),
        .\y[5] (_3560),
        .\y[6] (_3561),
        .\y[7] (_3562),
        .\y[8] (_3563),
        .\y[9] (_3564),
        .\y[10] (_3565),
        .\y[11] (_3566),
        .\y[12] (_3567),
        .\y[13] (_3568),
        .\y[14] (_3569),
        .\y[15] (_3570)
    );
    swap u51 (
        .\a[0] (_1540),
        .\a[1] (_1541),
        .\a[2] (_1542),
        .\a[3] (_1543),
        .\a[4] (_1544),
        .\a[5] (_1545),
        .\a[6] (_1546),
        .\a[7] (_1547),
        .\a[8] (_1548),
        .\a[9] (_1549),
        .\a[10] (_1550),
        .\a[11] (_1551),
        .\a[12] (_1552),
        .\a[13] (_1553),
        .\a[14] (_1554),
        .\a[15] (_1555),
        .\b[0] (_3279),
        .\b[1] (_3280),
        .\b[2] (_3281),
        .\b[3] (_3282),
        .\b[4] (_3283),
        .\b[5] (_3284),
        .\b[6] (_3285),
        .\b[7] (_3286),
        .\b[8] (_3287),
        .\b[9] (_3288),
        .\b[10] (_3289),
        .\b[11] (_3290),
        .\b[12] (_3291),
        .\b[13] (_3292),
        .\b[14] (_3293),
        .\b[15] (_3294),
        .\x[0] (_3604),
        .\x[1] (_3605),
        .\x[2] (_3606),
        .\x[3] (_3607),
        .\x[4] (_3608),
        .\x[5] (_3609),
        .\x[6] (_3610),
        .\x[7] (_3611),
        .\x[8] (_3612),
        .\x[9] (_3613),
        .\x[10] (_3614),
        .\x[11] (_3615),
        .\x[12] (_3616),
        .\x[13] (_3617),
        .\x[14] (_3618),
        .\x[15] (_3619),
        .\y[0] (_3620),
        .\y[1] (_3621),
        .\y[2] (_3622),
        .\y[3] (_3623),
        .\y[4] (_3624),
        .\y[5] (_3625),
        .\y[6] (_3626),
        .\y[7] (_3627),
        .\y[8] (_3628),
        .\y[9] (_3629),
        .\y[10] (_3630),
        .\y[11] (_3631),
        .\y[12] (_3632),
        .\y[13] (_3633),
        .\y[14] (_3634),
        .\y[15] (_3635)
    );
    swap u52 (
        .\a[0] (_1719),
        .\a[1] (_1720),
        .\a[2] (_1721),
        .\a[3] (_1722),
        .\a[4] (_1723),
        .\a[5] (_1724),
        .\a[6] (_1725),
        .\a[7] (_1726),
        .\a[8] (_1727),
        .\a[9] (_1728),
        .\a[10] (_1729),
        .\a[11] (_1730),
        .\a[12] (_1731),
        .\a[13] (_1732),
        .\a[14] (_1733),
        .\a[15] (_1734),
        .\b[0] (_3100),
        .\b[1] (_3101),
        .\b[2] (_3102),
        .\b[3] (_3103),
        .\b[4] (_3104),
        .\b[5] (_3105),
        .\b[6] (_3106),
        .\b[7] (_3107),
        .\b[8] (_3108),
        .\b[9] (_3109),
        .\b[10] (_3110),
        .\b[11] (_3111),
        .\b[12] (_3112),
        .\b[13] (_3113),
        .\b[14] (_3114),
        .\b[15] (_3115),
        .\x[0] (_3669),
        .\x[1] (_3670),
        .\x[2] (_3671),
        .\x[3] (_3672),
        .\x[4] (_3673),
        .\x[5] (_3674),
        .\x[6] (_3675),
        .\x[7] (_3676),
        .\x[8] (_3677),
        .\x[9] (_3678),
        .\x[10] (_3679),
        .\x[11] (_3680),
        .\x[12] (_3681),
        .\x[13] (_3682),
        .\x[14] (_3683),
        .\x[15] (_3684),
        .\y[0] (_3685),
        .\y[1] (_3686),
        .\y[2] (_3687),
        .\y[3] (_3688),
        .\y[4] (_3689),
        .\y[5] (_3690),
        .\y[6] (_3691),
        .\y[7] (_3692),
        .\y[8] (_3693),
        .\y[9] (_3694),
        .\y[10] (_3695),
        .\y[11] (_3696),
        .\y[12] (_3697),
        .\y[13] (_3698),
        .\y[14] (_3699),
        .\y[15] (_3700)
    );
    swap u53 (
        .\a[0] (_1735),
        .\a[1] (_1736),
        .\a[2] (_1737),
        .\a[3] (_1738),
        .\a[4] (_1739),
        .\a[5] (_1740),
        .\a[6] (_1741),
        .\a[7] (_1742),
        .\a[8] (_1743),
        .\a[9] (_1744),
        .\a[10] (_1745),
        .\a[11] (_1746),
        .\a[12] (_1747),
        .\a[13] (_1748),
        .\a[14] (_1749),
        .\a[15] (_1750),
        .\b[0] (_3084),
        .\b[1] (_3085),
        .\b[2] (_3086),
        .\b[3] (_3087),
        .\b[4] (_3088),
        .\b[5] (_3089),
        .\b[6] (_3090),
        .\b[7] (_3091),
        .\b[8] (_3092),
        .\b[9] (_3093),
        .\b[10] (_3094),
        .\b[11] (_3095),
        .\b[12] (_3096),
        .\b[13] (_3097),
        .\b[14] (_3098),
        .\b[15] (_3099),
        .\x[0] (_3734),
        .\x[1] (_3735),
        .\x[2] (_3736),
        .\x[3] (_3737),
        .\x[4] (_3738),
        .\x[5] (_3739),
        .\x[6] (_3740),
        .\x[7] (_3741),
        .\x[8] (_3742),
        .\x[9] (_3743),
        .\x[10] (_3744),
        .\x[11] (_3745),
        .\x[12] (_3746),
        .\x[13] (_3747),
        .\x[14] (_3748),
        .\x[15] (_3749),
        .\y[0] (_3750),
        .\y[1] (_3751),
        .\y[2] (_3752),
        .\y[3] (_3753),
        .\y[4] (_3754),
        .\y[5] (_3755),
        .\y[6] (_3756),
        .\y[7] (_3757),
        .\y[8] (_3758),
        .\y[9] (_3759),
        .\y[10] (_3760),
        .\y[11] (_3761),
        .\y[12] (_3762),
        .\y[13] (_3763),
        .\y[14] (_3764),
        .\y[15] (_3765)
    );
    swap u54 (
        .\a[0] (_1784),
        .\a[1] (_1785),
        .\a[2] (_1786),
        .\a[3] (_1787),
        .\a[4] (_1788),
        .\a[5] (_1789),
        .\a[6] (_1790),
        .\a[7] (_1791),
        .\a[8] (_1792),
        .\a[9] (_1793),
        .\a[10] (_1794),
        .\a[11] (_1795),
        .\a[12] (_1796),
        .\a[13] (_1797),
        .\a[14] (_1798),
        .\a[15] (_1799),
        .\b[0] (_3035),
        .\b[1] (_3036),
        .\b[2] (_3037),
        .\b[3] (_3038),
        .\b[4] (_3039),
        .\b[5] (_3040),
        .\b[6] (_3041),
        .\b[7] (_3042),
        .\b[8] (_3043),
        .\b[9] (_3044),
        .\b[10] (_3045),
        .\b[11] (_3046),
        .\b[12] (_3047),
        .\b[13] (_3048),
        .\b[14] (_3049),
        .\b[15] (_3050),
        .\x[0] (_3799),
        .\x[1] (_3800),
        .\x[2] (_3801),
        .\x[3] (_3802),
        .\x[4] (_3803),
        .\x[5] (_3804),
        .\x[6] (_3805),
        .\x[7] (_3806),
        .\x[8] (_3807),
        .\x[9] (_3808),
        .\x[10] (_3809),
        .\x[11] (_3810),
        .\x[12] (_3811),
        .\x[13] (_3812),
        .\x[14] (_3813),
        .\x[15] (_3814),
        .\y[0] (_3815),
        .\y[1] (_3816),
        .\y[2] (_3817),
        .\y[3] (_3818),
        .\y[4] (_3819),
        .\y[5] (_3820),
        .\y[6] (_3821),
        .\y[7] (_3822),
        .\y[8] (_3823),
        .\y[9] (_3824),
        .\y[10] (_3825),
        .\y[11] (_3826),
        .\y[12] (_3827),
        .\y[13] (_3828),
        .\y[14] (_3829),
        .\y[15] (_3830)
    );
    swap u55 (
        .\a[0] (_1800),
        .\a[1] (_1801),
        .\a[2] (_1802),
        .\a[3] (_1803),
        .\a[4] (_1804),
        .\a[5] (_1805),
        .\a[6] (_1806),
        .\a[7] (_1807),
        .\a[8] (_1808),
        .\a[9] (_1809),
        .\a[10] (_1810),
        .\a[11] (_1811),
        .\a[12] (_1812),
        .\a[13] (_1813),
        .\a[14] (_1814),
        .\a[15] (_1815),
        .\b[0] (_3019),
        .\b[1] (_3020),
        .\b[2] (_3021),
        .\b[3] (_3022),
        .\b[4] (_3023),
        .\b[5] (_3024),
        .\b[6] (_3025),
        .\b[7] (_3026),
        .\b[8] (_3027),
        .\b[9] (_3028),
        .\b[10] (_3029),
        .\b[11] (_3030),
        .\b[12] (_3031),
        .\b[13] (_3032),
        .\b[14] (_3033),
        .\b[15] (_3034),
        .\x[0] (_3864),
        .\x[1] (_3865),
        .\x[2] (_3866),
        .\x[3] (_3867),
        .\x[4] (_3868),
        .\x[5] (_3869),
        .\x[6] (_3870),
        .\x[7] (_3871),
        .\x[8] (_3872),
        .\x[9] (_3873),
        .\x[10] (_3874),
        .\x[11] (_3875),
        .\x[12] (_3876),
        .\x[13] (_3877),
        .\x[14] (_3878),
        .\x[15] (_3879),
        .\y[0] (_3880),
        .\y[1] (_3881),
        .\y[2] (_3882),
        .\y[3] (_3883),
        .\y[4] (_3884),
        .\y[5] (_3885),
        .\y[6] (_3886),
        .\y[7] (_3887),
        .\y[8] (_3888),
        .\y[9] (_3889),
        .\y[10] (_3890),
        .\y[11] (_3891),
        .\y[12] (_3892),
        .\y[13] (_3893),
        .\y[14] (_3894),
        .\y[15] (_3895)
    );
    swap u56 (
        .\a[0] (_3409),
        .\a[1] (_3410),
        .\a[2] (_3411),
        .\a[3] (_3412),
        .\a[4] (_3413),
        .\a[5] (_3414),
        .\a[6] (_3415),
        .\a[7] (_3416),
        .\a[8] (_3417),
        .\a[9] (_3418),
        .\a[10] (_3419),
        .\a[11] (_3420),
        .\a[12] (_3421),
        .\a[13] (_3422),
        .\a[14] (_3423),
        .\a[15] (_3424),
        .\b[0] (_3669),
        .\b[1] (_3670),
        .\b[2] (_3671),
        .\b[3] (_3672),
        .\b[4] (_3673),
        .\b[5] (_3674),
        .\b[6] (_3675),
        .\b[7] (_3676),
        .\b[8] (_3677),
        .\b[9] (_3678),
        .\b[10] (_3679),
        .\b[11] (_3680),
        .\b[12] (_3681),
        .\b[13] (_3682),
        .\b[14] (_3683),
        .\b[15] (_3684),
        .\x[0] (_3929),
        .\x[1] (_3930),
        .\x[2] (_3931),
        .\x[3] (_3932),
        .\x[4] (_3933),
        .\x[5] (_3934),
        .\x[6] (_3935),
        .\x[7] (_3936),
        .\x[8] (_3937),
        .\x[9] (_3938),
        .\x[10] (_3939),
        .\x[11] (_3940),
        .\x[12] (_3941),
        .\x[13] (_3942),
        .\x[14] (_3943),
        .\x[15] (_3944),
        .\y[0] (_3945),
        .\y[1] (_3946),
        .\y[2] (_3947),
        .\y[3] (_3948),
        .\y[4] (_3949),
        .\y[5] (_3950),
        .\y[6] (_3951),
        .\y[7] (_3952),
        .\y[8] (_3953),
        .\y[9] (_3954),
        .\y[10] (_3955),
        .\y[11] (_3956),
        .\y[12] (_3957),
        .\y[13] (_3958),
        .\y[14] (_3959),
        .\y[15] (_3960)
    );
    swap u57 (
        .\a[0] (_3474),
        .\a[1] (_3475),
        .\a[2] (_3476),
        .\a[3] (_3477),
        .\a[4] (_3478),
        .\a[5] (_3479),
        .\a[6] (_3480),
        .\a[7] (_3481),
        .\a[8] (_3482),
        .\a[9] (_3483),
        .\a[10] (_3484),
        .\a[11] (_3485),
        .\a[12] (_3486),
        .\a[13] (_3487),
        .\a[14] (_3488),
        .\a[15] (_3489),
        .\b[0] (_3734),
        .\b[1] (_3735),
        .\b[2] (_3736),
        .\b[3] (_3737),
        .\b[4] (_3738),
        .\b[5] (_3739),
        .\b[6] (_3740),
        .\b[7] (_3741),
        .\b[8] (_3742),
        .\b[9] (_3743),
        .\b[10] (_3744),
        .\b[11] (_3745),
        .\b[12] (_3746),
        .\b[13] (_3747),
        .\b[14] (_3748),
        .\b[15] (_3749),
        .\x[0] (_3994),
        .\x[1] (_3995),
        .\x[2] (_3996),
        .\x[3] (_3997),
        .\x[4] (_3998),
        .\x[5] (_3999),
        .\x[6] (_4000),
        .\x[7] (_4001),
        .\x[8] (_4002),
        .\x[9] (_4003),
        .\x[10] (_4004),
        .\x[11] (_4005),
        .\x[12] (_4006),
        .\x[13] (_4007),
        .\x[14] (_4008),
        .\x[15] (_4009),
        .\y[0] (_4010),
        .\y[1] (_4011),
        .\y[2] (_4012),
        .\y[3] (_4013),
        .\y[4] (_4014),
        .\y[5] (_4015),
        .\y[6] (_4016),
        .\y[7] (_4017),
        .\y[8] (_4018),
        .\y[9] (_4019),
        .\y[10] (_4020),
        .\y[11] (_4021),
        .\y[12] (_4022),
        .\y[13] (_4023),
        .\y[14] (_4024),
        .\y[15] (_4025)
    );
    swap u58 (
        .\a[0] (_3539),
        .\a[1] (_3540),
        .\a[2] (_3541),
        .\a[3] (_3542),
        .\a[4] (_3543),
        .\a[5] (_3544),
        .\a[6] (_3545),
        .\a[7] (_3546),
        .\a[8] (_3547),
        .\a[9] (_3548),
        .\a[10] (_3549),
        .\a[11] (_3550),
        .\a[12] (_3551),
        .\a[13] (_3552),
        .\a[14] (_3553),
        .\a[15] (_3554),
        .\b[0] (_3799),
        .\b[1] (_3800),
        .\b[2] (_3801),
        .\b[3] (_3802),
        .\b[4] (_3803),
        .\b[5] (_3804),
        .\b[6] (_3805),
        .\b[7] (_3806),
        .\b[8] (_3807),
        .\b[9] (_3808),
        .\b[10] (_3809),
        .\b[11] (_3810),
        .\b[12] (_3811),
        .\b[13] (_3812),
        .\b[14] (_3813),
        .\b[15] (_3814),
        .\x[0] (_4059),
        .\x[1] (_4060),
        .\x[2] (_4061),
        .\x[3] (_4062),
        .\x[4] (_4063),
        .\x[5] (_4064),
        .\x[6] (_4065),
        .\x[7] (_4066),
        .\x[8] (_4067),
        .\x[9] (_4068),
        .\x[10] (_4069),
        .\x[11] (_4070),
        .\x[12] (_4071),
        .\x[13] (_4072),
        .\x[14] (_4073),
        .\x[15] (_4074),
        .\y[0] (_4075),
        .\y[1] (_4076),
        .\y[2] (_4077),
        .\y[3] (_4078),
        .\y[4] (_4079),
        .\y[5] (_4080),
        .\y[6] (_4081),
        .\y[7] (_4082),
        .\y[8] (_4083),
        .\y[9] (_4084),
        .\y[10] (_4085),
        .\y[11] (_4086),
        .\y[12] (_4087),
        .\y[13] (_4088),
        .\y[14] (_4089),
        .\y[15] (_4090)
    );
    swap u59 (
        .\a[0] (_3604),
        .\a[1] (_3605),
        .\a[2] (_3606),
        .\a[3] (_3607),
        .\a[4] (_3608),
        .\a[5] (_3609),
        .\a[6] (_3610),
        .\a[7] (_3611),
        .\a[8] (_3612),
        .\a[9] (_3613),
        .\a[10] (_3614),
        .\a[11] (_3615),
        .\a[12] (_3616),
        .\a[13] (_3617),
        .\a[14] (_3618),
        .\a[15] (_3619),
        .\b[0] (_3864),
        .\b[1] (_3865),
        .\b[2] (_3866),
        .\b[3] (_3867),
        .\b[4] (_3868),
        .\b[5] (_3869),
        .\b[6] (_3870),
        .\b[7] (_3871),
        .\b[8] (_3872),
        .\b[9] (_3873),
        .\b[10] (_3874),
        .\b[11] (_3875),
        .\b[12] (_3876),
        .\b[13] (_3877),
        .\b[14] (_3878),
        .\b[15] (_3879),
        .\x[0] (_4124),
        .\x[1] (_4125),
        .\x[2] (_4126),
        .\x[3] (_4127),
        .\x[4] (_4128),
        .\x[5] (_4129),
        .\x[6] (_4130),
        .\x[7] (_4131),
        .\x[8] (_4132),
        .\x[9] (_4133),
        .\x[10] (_4134),
        .\x[11] (_4135),
        .\x[12] (_4136),
        .\x[13] (_4137),
        .\x[14] (_4138),
        .\x[15] (_4139),
        .\y[0] (_4140),
        .\y[1] (_4141),
        .\y[2] (_4142),
        .\y[3] (_4143),
        .\y[4] (_4144),
        .\y[5] (_4145),
        .\y[6] (_4146),
        .\y[7] (_4147),
        .\y[8] (_4148),
        .\y[9] (_4149),
        .\y[10] (_4150),
        .\y[11] (_4151),
        .\y[12] (_4152),
        .\y[13] (_4153),
        .\y[14] (_4154),
        .\y[15] (_4155)
    );
    swap u60 (
        .\a[0] (_3929),
        .\a[1] (_3930),
        .\a[2] (_3931),
        .\a[3] (_3932),
        .\a[4] (_3933),
        .\a[5] (_3934),
        .\a[6] (_3935),
        .\a[7] (_3936),
        .\a[8] (_3937),
        .\a[9] (_3938),
        .\a[10] (_3939),
        .\a[11] (_3940),
        .\a[12] (_3941),
        .\a[13] (_3942),
        .\a[14] (_3943),
        .\a[15] (_3944),
        .\b[0] (_4059),
        .\b[1] (_4060),
        .\b[2] (_4061),
        .\b[3] (_4062),
        .\b[4] (_4063),
        .\b[5] (_4064),
        .\b[6] (_4065),
        .\b[7] (_4066),
        .\b[8] (_4067),
        .\b[9] (_4068),
        .\b[10] (_4069),
        .\b[11] (_4070),
        .\b[12] (_4071),
        .\b[13] (_4072),
        .\b[14] (_4073),
        .\b[15] (_4074),
        .\x[0] (_4189),
        .\x[1] (_4190),
        .\x[2] (_4191),
        .\x[3] (_4192),
        .\x[4] (_4193),
        .\x[5] (_4194),
        .\x[6] (_4195),
        .\x[7] (_4196),
        .\x[8] (_4197),
        .\x[9] (_4198),
        .\x[10] (_4199),
        .\x[11] (_4200),
        .\x[12] (_4201),
        .\x[13] (_4202),
        .\x[14] (_4203),
        .\x[15] (_4204),
        .\y[0] (_4205),
        .\y[1] (_4206),
        .\y[2] (_4207),
        .\y[3] (_4208),
        .\y[4] (_4209),
        .\y[5] (_4210),
        .\y[6] (_4211),
        .\y[7] (_4212),
        .\y[8] (_4213),
        .\y[9] (_4214),
        .\y[10] (_4215),
        .\y[11] (_4216),
        .\y[12] (_4217),
        .\y[13] (_4218),
        .\y[14] (_4219),
        .\y[15] (_4220)
    );
    swap u61 (
        .\a[0] (_3994),
        .\a[1] (_3995),
        .\a[2] (_3996),
        .\a[3] (_3997),
        .\a[4] (_3998),
        .\a[5] (_3999),
        .\a[6] (_4000),
        .\a[7] (_4001),
        .\a[8] (_4002),
        .\a[9] (_4003),
        .\a[10] (_4004),
        .\a[11] (_4005),
        .\a[12] (_4006),
        .\a[13] (_4007),
        .\a[14] (_4008),
        .\a[15] (_4009),
        .\b[0] (_4124),
        .\b[1] (_4125),
        .\b[2] (_4126),
        .\b[3] (_4127),
        .\b[4] (_4128),
        .\b[5] (_4129),
        .\b[6] (_4130),
        .\b[7] (_4131),
        .\b[8] (_4132),
        .\b[9] (_4133),
        .\b[10] (_4134),
        .\b[11] (_4135),
        .\b[12] (_4136),
        .\b[13] (_4137),
        .\b[14] (_4138),
        .\b[15] (_4139),
        .\x[0] (_4254),
        .\x[1] (_4255),
        .\x[2] (_4256),
        .\x[3] (_4257),
        .\x[4] (_4258),
        .\x[5] (_4259),
        .\x[6] (_4260),
        .\x[7] (_4261),
        .\x[8] (_4262),
        .\x[9] (_4263),
        .\x[10] (_4264),
        .\x[11] (_4265),
        .\x[12] (_4266),
        .\x[13] (_4267),
        .\x[14] (_4268),
        .\x[15] (_4269),
        .\y[0] (_4270),
        .\y[1] (_4271),
        .\y[2] (_4272),
        .\y[3] (_4273),
        .\y[4] (_4274),
        .\y[5] (_4275),
        .\y[6] (_4276),
        .\y[7] (_4277),
        .\y[8] (_4278),
        .\y[9] (_4279),
        .\y[10] (_4280),
        .\y[11] (_4281),
        .\y[12] (_4282),
        .\y[13] (_4283),
        .\y[14] (_4284),
        .\y[15] (_4285)
    );
    swap u62 (
        .\a[0] (_4189),
        .\a[1] (_4190),
        .\a[2] (_4191),
        .\a[3] (_4192),
        .\a[4] (_4193),
        .\a[5] (_4194),
        .\a[6] (_4195),
        .\a[7] (_4196),
        .\a[8] (_4197),
        .\a[9] (_4198),
        .\a[10] (_4199),
        .\a[11] (_4200),
        .\a[12] (_4201),
        .\a[13] (_4202),
        .\a[14] (_4203),
        .\a[15] (_4204),
        .\b[0] (_4254),
        .\b[1] (_4255),
        .\b[2] (_4256),
        .\b[3] (_4257),
        .\b[4] (_4258),
        .\b[5] (_4259),
        .\b[6] (_4260),
        .\b[7] (_4261),
        .\b[8] (_4262),
        .\b[9] (_4263),
        .\b[10] (_4264),
        .\b[11] (_4265),
        .\b[12] (_4266),
        .\b[13] (_4267),
        .\b[14] (_4268),
        .\b[15] (_4269),
        .\x[0] (_4319),
        .\x[1] (_4320),
        .\x[2] (_4321),
        .\x[3] (_4322),
        .\x[4] (_4323),
        .\x[5] (_4324),
        .\x[6] (_4325),
        .\x[7] (_4326),
        .\x[8] (_4327),
        .\x[9] (_4328),
        .\x[10] (_4329),
        .\x[11] (_4330),
        .\x[12] (_4331),
        .\x[13] (_4332),
        .\x[14] (_4333),
        .\x[15] (_4334),
        .\y[0] (_4335),
        .\y[1] (_4336),
        .\y[2] (_4337),
        .\y[3] (_4338),
        .\y[4] (_4339),
        .\y[5] (_4340),
        .\y[6] (_4341),
        .\y[7] (_4342),
        .\y[8] (_4343),
        .\y[9] (_4344),
        .\y[10] (_4345),
        .\y[11] (_4346),
        .\y[12] (_4347),
        .\y[13] (_4348),
        .\y[14] (_4349),
        .\y[15] (_4350)
    );
    swap u63 (
        .\a[0] (_4205),
        .\a[1] (_4206),
        .\a[2] (_4207),
        .\a[3] (_4208),
        .\a[4] (_4209),
        .\a[5] (_4210),
        .\a[6] (_4211),
        .\a[7] (_4212),
        .\a[8] (_4213),
        .\a[9] (_4214),
        .\a[10] (_4215),
        .\a[11] (_4216),
        .\a[12] (_4217),
        .\a[13] (_4218),
        .\a[14] (_4219),
        .\a[15] (_4220),
        .\b[0] (_4270),
        .\b[1] (_4271),
        .\b[2] (_4272),
        .\b[3] (_4273),
        .\b[4] (_4274),
        .\b[5] (_4275),
        .\b[6] (_4276),
        .\b[7] (_4277),
        .\b[8] (_4278),
        .\b[9] (_4279),
        .\b[10] (_4280),
        .\b[11] (_4281),
        .\b[12] (_4282),
        .\b[13] (_4283),
        .\b[14] (_4284),
        .\b[15] (_4285),
        .\x[0] (_4384),
        .\x[1] (_4385),
        .\x[2] (_4386),
        .\x[3] (_4387),
        .\x[4] (_4388),
        .\x[5] (_4389),
        .\x[6] (_4390),
        .\x[7] (_4391),
        .\x[8] (_4392),
        .\x[9] (_4393),
        .\x[10] (_4394),
        .\x[11] (_4395),
        .\x[12] (_4396),
        .\x[13] (_4397),
        .\x[14] (_4398),
        .\x[15] (_4399),
        .\y[0] (_4400),
        .\y[1] (_4401),
        .\y[2] (_4402),
        .\y[3] (_4403),
        .\y[4] (_4404),
        .\y[5] (_4405),
        .\y[6] (_4406),
        .\y[7] (_4407),
        .\y[8] (_4408),
        .\y[9] (_4409),
        .\y[10] (_4410),
        .\y[11] (_4411),
        .\y[12] (_4412),
        .\y[13] (_4413),
        .\y[14] (_4414),
        .\y[15] (_4415)
    );
    swap u64 (
        .\a[0] (_3945),
        .\a[1] (_3946),
        .\a[2] (_3947),
        .\a[3] (_3948),
        .\a[4] (_3949),
        .\a[5] (_3950),
        .\a[6] (_3951),
        .\a[7] (_3952),
        .\a[8] (_3953),
        .\a[9] (_3954),
        .\a[10] (_3955),
        .\a[11] (_3956),
        .\a[12] (_3957),
        .\a[13] (_3958),
        .\a[14] (_3959),
        .\a[15] (_3960),
        .\b[0] (_4075),
        .\b[1] (_4076),
        .\b[2] (_4077),
        .\b[3] (_4078),
        .\b[4] (_4079),
        .\b[5] (_4080),
        .\b[6] (_4081),
        .\b[7] (_4082),
        .\b[8] (_4083),
        .\b[9] (_4084),
        .\b[10] (_4085),
        .\b[11] (_4086),
        .\b[12] (_4087),
        .\b[13] (_4088),
        .\b[14] (_4089),
        .\b[15] (_4090),
        .\x[0] (_4449),
        .\x[1] (_4450),
        .\x[2] (_4451),
        .\x[3] (_4452),
        .\x[4] (_4453),
        .\x[5] (_4454),
        .\x[6] (_4455),
        .\x[7] (_4456),
        .\x[8] (_4457),
        .\x[9] (_4458),
        .\x[10] (_4459),
        .\x[11] (_4460),
        .\x[12] (_4461),
        .\x[13] (_4462),
        .\x[14] (_4463),
        .\x[15] (_4464),
        .\y[0] (_4465),
        .\y[1] (_4466),
        .\y[2] (_4467),
        .\y[3] (_4468),
        .\y[4] (_4469),
        .\y[5] (_4470),
        .\y[6] (_4471),
        .\y[7] (_4472),
        .\y[8] (_4473),
        .\y[9] (_4474),
        .\y[10] (_4475),
        .\y[11] (_4476),
        .\y[12] (_4477),
        .\y[13] (_4478),
        .\y[14] (_4479),
        .\y[15] (_4480)
    );
    swap u65 (
        .\a[0] (_4010),
        .\a[1] (_4011),
        .\a[2] (_4012),
        .\a[3] (_4013),
        .\a[4] (_4014),
        .\a[5] (_4015),
        .\a[6] (_4016),
        .\a[7] (_4017),
        .\a[8] (_4018),
        .\a[9] (_4019),
        .\a[10] (_4020),
        .\a[11] (_4021),
        .\a[12] (_4022),
        .\a[13] (_4023),
        .\a[14] (_4024),
        .\a[15] (_4025),
        .\b[0] (_4140),
        .\b[1] (_4141),
        .\b[2] (_4142),
        .\b[3] (_4143),
        .\b[4] (_4144),
        .\b[5] (_4145),
        .\b[6] (_4146),
        .\b[7] (_4147),
        .\b[8] (_4148),
        .\b[9] (_4149),
        .\b[10] (_4150),
        .\b[11] (_4151),
        .\b[12] (_4152),
        .\b[13] (_4153),
        .\b[14] (_4154),
        .\b[15] (_4155),
        .\x[0] (_4514),
        .\x[1] (_4515),
        .\x[2] (_4516),
        .\x[3] (_4517),
        .\x[4] (_4518),
        .\x[5] (_4519),
        .\x[6] (_4520),
        .\x[7] (_4521),
        .\x[8] (_4522),
        .\x[9] (_4523),
        .\x[10] (_4524),
        .\x[11] (_4525),
        .\x[12] (_4526),
        .\x[13] (_4527),
        .\x[14] (_4528),
        .\x[15] (_4529),
        .\y[0] (_4530),
        .\y[1] (_4531),
        .\y[2] (_4532),
        .\y[3] (_4533),
        .\y[4] (_4534),
        .\y[5] (_4535),
        .\y[6] (_4536),
        .\y[7] (_4537),
        .\y[8] (_4538),
        .\y[9] (_4539),
        .\y[10] (_4540),
        .\y[11] (_4541),
        .\y[12] (_4542),
        .\y[13] (_4543),
        .\y[14] (_4544),
        .\y[15] (_4545)
    );
    swap u66 (
        .\a[0] (_4449),
        .\a[1] (_4450),
        .\a[2] (_4451),
        .\a[3] (_4452),
        .\a[4] (_4453),
        .\a[5] (_4454),
        .\a[6] (_4455),
        .\a[7] (_4456),
        .\a[8] (_4457),
        .\a[9] (_4458),
        .\a[10] (_4459),
        .\a[11] (_4460),
        .\a[12] (_4461),
        .\a[13] (_4462),
        .\a[14] (_4463),
        .\a[15] (_4464),
        .\b[0] (_4514),
        .\b[1] (_4515),
        .\b[2] (_4516),
        .\b[3] (_4517),
        .\b[4] (_4518),
        .\b[5] (_4519),
        .\b[6] (_4520),
        .\b[7] (_4521),
        .\b[8] (_4522),
        .\b[9] (_4523),
        .\b[10] (_4524),
        .\b[11] (_4525),
        .\b[12] (_4526),
        .\b[13] (_4527),
        .\b[14] (_4528),
        .\b[15] (_4529),
        .\x[0] (_4579),
        .\x[1] (_4580),
        .\x[2] (_4581),
        .\x[3] (_4582),
        .\x[4] (_4583),
        .\x[5] (_4584),
        .\x[6] (_4585),
        .\x[7] (_4586),
        .\x[8] (_4587),
        .\x[9] (_4588),
        .\x[10] (_4589),
        .\x[11] (_4590),
        .\x[12] (_4591),
        .\x[13] (_4592),
        .\x[14] (_4593),
        .\x[15] (_4594),
        .\y[0] (_4595),
        .\y[1] (_4596),
        .\y[2] (_4597),
        .\y[3] (_4598),
        .\y[4] (_4599),
        .\y[5] (_4600),
        .\y[6] (_4601),
        .\y[7] (_4602),
        .\y[8] (_4603),
        .\y[9] (_4604),
        .\y[10] (_4605),
        .\y[11] (_4606),
        .\y[12] (_4607),
        .\y[13] (_4608),
        .\y[14] (_4609),
        .\y[15] (_4610)
    );
    swap u67 (
        .\a[0] (_4465),
        .\a[1] (_4466),
        .\a[2] (_4467),
        .\a[3] (_4468),
        .\a[4] (_4469),
        .\a[5] (_4470),
        .\a[6] (_4471),
        .\a[7] (_4472),
        .\a[8] (_4473),
        .\a[9] (_4474),
        .\a[10] (_4475),
        .\a[11] (_4476),
        .\a[12] (_4477),
        .\a[13] (_4478),
        .\a[14] (_4479),
        .\a[15] (_4480),
        .\b[0] (_4530),
        .\b[1] (_4531),
        .\b[2] (_4532),
        .\b[3] (_4533),
        .\b[4] (_4534),
        .\b[5] (_4535),
        .\b[6] (_4536),
        .\b[7] (_4537),
        .\b[8] (_4538),
        .\b[9] (_4539),
        .\b[10] (_4540),
        .\b[11] (_4541),
        .\b[12] (_4542),
        .\b[13] (_4543),
        .\b[14] (_4544),
        .\b[15] (_4545),
        .\x[0] (_4644),
        .\x[1] (_4645),
        .\x[2] (_4646),
        .\x[3] (_4647),
        .\x[4] (_4648),
        .\x[5] (_4649),
        .\x[6] (_4650),
        .\x[7] (_4651),
        .\x[8] (_4652),
        .\x[9] (_4653),
        .\x[10] (_4654),
        .\x[11] (_4655),
        .\x[12] (_4656),
        .\x[13] (_4657),
        .\x[14] (_4658),
        .\x[15] (_4659),
        .\y[0] (_4660),
        .\y[1] (_4661),
        .\y[2] (_4662),
        .\y[3] (_4663),
        .\y[4] (_4664),
        .\y[5] (_4665),
        .\y[6] (_4666),
        .\y[7] (_4667),
        .\y[8] (_4668),
        .\y[9] (_4669),
        .\y[10] (_4670),
        .\y[11] (_4671),
        .\y[12] (_4672),
        .\y[13] (_4673),
        .\y[14] (_4674),
        .\y[15] (_4675)
    );
    swap u68 (
        .\a[0] (_3425),
        .\a[1] (_3426),
        .\a[2] (_3427),
        .\a[3] (_3428),
        .\a[4] (_3429),
        .\a[5] (_3430),
        .\a[6] (_3431),
        .\a[7] (_3432),
        .\a[8] (_3433),
        .\a[9] (_3434),
        .\a[10] (_3435),
        .\a[11] (_3436),
        .\a[12] (_3437),
        .\a[13] (_3438),
        .\a[14] (_3439),
        .\a[15] (_3440),
        .\b[0] (_3685),
        .\b[1] (_3686),
        .\b[2] (_3687),
        .\b[3] (_3688),
        .\b[4] (_3689),
        .\b[5] (_3690),
        .\b[6] (_3691),
        .\b[7] (_3692),
        .\b[8] (_3693),
        .\b[9] (_3694),
        .\b[10] (_3695),
        .\b[11] (_3696),
        .\b[12] (_3697),
        .\b[13] (_3698),
        .\b[14] (_3699),
        .\b[15] (_3700),
        .\x[0] (_4709),
        .\x[1] (_4710),
        .\x[2] (_4711),
        .\x[3] (_4712),
        .\x[4] (_4713),
        .\x[5] (_4714),
        .\x[6] (_4715),
        .\x[7] (_4716),
        .\x[8] (_4717),
        .\x[9] (_4718),
        .\x[10] (_4719),
        .\x[11] (_4720),
        .\x[12] (_4721),
        .\x[13] (_4722),
        .\x[14] (_4723),
        .\x[15] (_4724),
        .\y[0] (_4725),
        .\y[1] (_4726),
        .\y[2] (_4727),
        .\y[3] (_4728),
        .\y[4] (_4729),
        .\y[5] (_4730),
        .\y[6] (_4731),
        .\y[7] (_4732),
        .\y[8] (_4733),
        .\y[9] (_4734),
        .\y[10] (_4735),
        .\y[11] (_4736),
        .\y[12] (_4737),
        .\y[13] (_4738),
        .\y[14] (_4739),
        .\y[15] (_4740)
    );
    swap u69 (
        .\a[0] (_3490),
        .\a[1] (_3491),
        .\a[2] (_3492),
        .\a[3] (_3493),
        .\a[4] (_3494),
        .\a[5] (_3495),
        .\a[6] (_3496),
        .\a[7] (_3497),
        .\a[8] (_3498),
        .\a[9] (_3499),
        .\a[10] (_3500),
        .\a[11] (_3501),
        .\a[12] (_3502),
        .\a[13] (_3503),
        .\a[14] (_3504),
        .\a[15] (_3505),
        .\b[0] (_3750),
        .\b[1] (_3751),
        .\b[2] (_3752),
        .\b[3] (_3753),
        .\b[4] (_3754),
        .\b[5] (_3755),
        .\b[6] (_3756),
        .\b[7] (_3757),
        .\b[8] (_3758),
        .\b[9] (_3759),
        .\b[10] (_3760),
        .\b[11] (_3761),
        .\b[12] (_3762),
        .\b[13] (_3763),
        .\b[14] (_3764),
        .\b[15] (_3765),
        .\x[0] (_4774),
        .\x[1] (_4775),
        .\x[2] (_4776),
        .\x[3] (_4777),
        .\x[4] (_4778),
        .\x[5] (_4779),
        .\x[6] (_4780),
        .\x[7] (_4781),
        .\x[8] (_4782),
        .\x[9] (_4783),
        .\x[10] (_4784),
        .\x[11] (_4785),
        .\x[12] (_4786),
        .\x[13] (_4787),
        .\x[14] (_4788),
        .\x[15] (_4789),
        .\y[0] (_4790),
        .\y[1] (_4791),
        .\y[2] (_4792),
        .\y[3] (_4793),
        .\y[4] (_4794),
        .\y[5] (_4795),
        .\y[6] (_4796),
        .\y[7] (_4797),
        .\y[8] (_4798),
        .\y[9] (_4799),
        .\y[10] (_4800),
        .\y[11] (_4801),
        .\y[12] (_4802),
        .\y[13] (_4803),
        .\y[14] (_4804),
        .\y[15] (_4805)
    );
    swap u70 (
        .\a[0] (_3555),
        .\a[1] (_3556),
        .\a[2] (_3557),
        .\a[3] (_3558),
        .\a[4] (_3559),
        .\a[5] (_3560),
        .\a[6] (_3561),
        .\a[7] (_3562),
        .\a[8] (_3563),
        .\a[9] (_3564),
        .\a[10] (_3565),
        .\a[11] (_3566),
        .\a[12] (_3567),
        .\a[13] (_3568),
        .\a[14] (_3569),
        .\a[15] (_3570),
        .\b[0] (_3815),
        .\b[1] (_3816),
        .\b[2] (_3817),
        .\b[3] (_3818),
        .\b[4] (_3819),
        .\b[5] (_3820),
        .\b[6] (_3821),
        .\b[7] (_3822),
        .\b[8] (_3823),
        .\b[9] (_3824),
        .\b[10] (_3825),
        .\b[11] (_3826),
        .\b[12] (_3827),
        .\b[13] (_3828),
        .\b[14] (_3829),
        .\b[15] (_3830),
        .\x[0] (_4839),
        .\x[1] (_4840),
        .\x[2] (_4841),
        .\x[3] (_4842),
        .\x[4] (_4843),
        .\x[5] (_4844),
        .\x[6] (_4845),
        .\x[7] (_4846),
        .\x[8] (_4847),
        .\x[9] (_4848),
        .\x[10] (_4849),
        .\x[11] (_4850),
        .\x[12] (_4851),
        .\x[13] (_4852),
        .\x[14] (_4853),
        .\x[15] (_4854),
        .\y[0] (_4855),
        .\y[1] (_4856),
        .\y[2] (_4857),
        .\y[3] (_4858),
        .\y[4] (_4859),
        .\y[5] (_4860),
        .\y[6] (_4861),
        .\y[7] (_4862),
        .\y[8] (_4863),
        .\y[9] (_4864),
        .\y[10] (_4865),
        .\y[11] (_4866),
        .\y[12] (_4867),
        .\y[13] (_4868),
        .\y[14] (_4869),
        .\y[15] (_4870)
    );
    swap u71 (
        .\a[0] (_3620),
        .\a[1] (_3621),
        .\a[2] (_3622),
        .\a[3] (_3623),
        .\a[4] (_3624),
        .\a[5] (_3625),
        .\a[6] (_3626),
        .\a[7] (_3627),
        .\a[8] (_3628),
        .\a[9] (_3629),
        .\a[10] (_3630),
        .\a[11] (_3631),
        .\a[12] (_3632),
        .\a[13] (_3633),
        .\a[14] (_3634),
        .\a[15] (_3635),
        .\b[0] (_3880),
        .\b[1] (_3881),
        .\b[2] (_3882),
        .\b[3] (_3883),
        .\b[4] (_3884),
        .\b[5] (_3885),
        .\b[6] (_3886),
        .\b[7] (_3887),
        .\b[8] (_3888),
        .\b[9] (_3889),
        .\b[10] (_3890),
        .\b[11] (_3891),
        .\b[12] (_3892),
        .\b[13] (_3893),
        .\b[14] (_3894),
        .\b[15] (_3895),
        .\x[0] (_4904),
        .\x[1] (_4905),
        .\x[2] (_4906),
        .\x[3] (_4907),
        .\x[4] (_4908),
        .\x[5] (_4909),
        .\x[6] (_4910),
        .\x[7] (_4911),
        .\x[8] (_4912),
        .\x[9] (_4913),
        .\x[10] (_4914),
        .\x[11] (_4915),
        .\x[12] (_4916),
        .\x[13] (_4917),
        .\x[14] (_4918),
        .\x[15] (_4919),
        .\y[0] (_4920),
        .\y[1] (_4921),
        .\y[2] (_4922),
        .\y[3] (_4923),
        .\y[4] (_4924),
        .\y[5] (_4925),
        .\y[6] (_4926),
        .\y[7] (_4927),
        .\y[8] (_4928),
        .\y[9] (_4929),
        .\y[10] (_4930),
        .\y[11] (_4931),
        .\y[12] (_4932),
        .\y[13] (_4933),
        .\y[14] (_4934),
        .\y[15] (_4935)
    );
    swap u72 (
        .\a[0] (_4709),
        .\a[1] (_4710),
        .\a[2] (_4711),
        .\a[3] (_4712),
        .\a[4] (_4713),
        .\a[5] (_4714),
        .\a[6] (_4715),
        .\a[7] (_4716),
        .\a[8] (_4717),
        .\a[9] (_4718),
        .\a[10] (_4719),
        .\a[11] (_4720),
        .\a[12] (_4721),
        .\a[13] (_4722),
        .\a[14] (_4723),
        .\a[15] (_4724),
        .\b[0] (_4839),
        .\b[1] (_4840),
        .\b[2] (_4841),
        .\b[3] (_4842),
        .\b[4] (_4843),
        .\b[5] (_4844),
        .\b[6] (_4845),
        .\b[7] (_4846),
        .\b[8] (_4847),
        .\b[9] (_4848),
        .\b[10] (_4849),
        .\b[11] (_4850),
        .\b[12] (_4851),
        .\b[13] (_4852),
        .\b[14] (_4853),
        .\b[15] (_4854),
        .\x[0] (_4969),
        .\x[1] (_4970),
        .\x[2] (_4971),
        .\x[3] (_4972),
        .\x[4] (_4973),
        .\x[5] (_4974),
        .\x[6] (_4975),
        .\x[7] (_4976),
        .\x[8] (_4977),
        .\x[9] (_4978),
        .\x[10] (_4979),
        .\x[11] (_4980),
        .\x[12] (_4981),
        .\x[13] (_4982),
        .\x[14] (_4983),
        .\x[15] (_4984),
        .\y[0] (_4985),
        .\y[1] (_4986),
        .\y[2] (_4987),
        .\y[3] (_4988),
        .\y[4] (_4989),
        .\y[5] (_4990),
        .\y[6] (_4991),
        .\y[7] (_4992),
        .\y[8] (_4993),
        .\y[9] (_4994),
        .\y[10] (_4995),
        .\y[11] (_4996),
        .\y[12] (_4997),
        .\y[13] (_4998),
        .\y[14] (_4999),
        .\y[15] (_5000)
    );
    swap u73 (
        .\a[0] (_4774),
        .\a[1] (_4775),
        .\a[2] (_4776),
        .\a[3] (_4777),
        .\a[4] (_4778),
        .\a[5] (_4779),
        .\a[6] (_4780),
        .\a[7] (_4781),
        .\a[8] (_4782),
        .\a[9] (_4783),
        .\a[10] (_4784),
        .\a[11] (_4785),
        .\a[12] (_4786),
        .\a[13] (_4787),
        .\a[14] (_4788),
        .\a[15] (_4789),
        .\b[0] (_4904),
        .\b[1] (_4905),
        .\b[2] (_4906),
        .\b[3] (_4907),
        .\b[4] (_4908),
        .\b[5] (_4909),
        .\b[6] (_4910),
        .\b[7] (_4911),
        .\b[8] (_4912),
        .\b[9] (_4913),
        .\b[10] (_4914),
        .\b[11] (_4915),
        .\b[12] (_4916),
        .\b[13] (_4917),
        .\b[14] (_4918),
        .\b[15] (_4919),
        .\x[0] (_5034),
        .\x[1] (_5035),
        .\x[2] (_5036),
        .\x[3] (_5037),
        .\x[4] (_5038),
        .\x[5] (_5039),
        .\x[6] (_5040),
        .\x[7] (_5041),
        .\x[8] (_5042),
        .\x[9] (_5043),
        .\x[10] (_5044),
        .\x[11] (_5045),
        .\x[12] (_5046),
        .\x[13] (_5047),
        .\x[14] (_5048),
        .\x[15] (_5049),
        .\y[0] (_5050),
        .\y[1] (_5051),
        .\y[2] (_5052),
        .\y[3] (_5053),
        .\y[4] (_5054),
        .\y[5] (_5055),
        .\y[6] (_5056),
        .\y[7] (_5057),
        .\y[8] (_5058),
        .\y[9] (_5059),
        .\y[10] (_5060),
        .\y[11] (_5061),
        .\y[12] (_5062),
        .\y[13] (_5063),
        .\y[14] (_5064),
        .\y[15] (_5065)
    );
    swap u74 (
        .\a[0] (_4969),
        .\a[1] (_4970),
        .\a[2] (_4971),
        .\a[3] (_4972),
        .\a[4] (_4973),
        .\a[5] (_4974),
        .\a[6] (_4975),
        .\a[7] (_4976),
        .\a[8] (_4977),
        .\a[9] (_4978),
        .\a[10] (_4979),
        .\a[11] (_4980),
        .\a[12] (_4981),
        .\a[13] (_4982),
        .\a[14] (_4983),
        .\a[15] (_4984),
        .\b[0] (_5034),
        .\b[1] (_5035),
        .\b[2] (_5036),
        .\b[3] (_5037),
        .\b[4] (_5038),
        .\b[5] (_5039),
        .\b[6] (_5040),
        .\b[7] (_5041),
        .\b[8] (_5042),
        .\b[9] (_5043),
        .\b[10] (_5044),
        .\b[11] (_5045),
        .\b[12] (_5046),
        .\b[13] (_5047),
        .\b[14] (_5048),
        .\b[15] (_5049),
        .\x[0] (_5099),
        .\x[1] (_5100),
        .\x[2] (_5101),
        .\x[3] (_5102),
        .\x[4] (_5103),
        .\x[5] (_5104),
        .\x[6] (_5105),
        .\x[7] (_5106),
        .\x[8] (_5107),
        .\x[9] (_5108),
        .\x[10] (_5109),
        .\x[11] (_5110),
        .\x[12] (_5111),
        .\x[13] (_5112),
        .\x[14] (_5113),
        .\x[15] (_5114),
        .\y[0] (_5115),
        .\y[1] (_5116),
        .\y[2] (_5117),
        .\y[3] (_5118),
        .\y[4] (_5119),
        .\y[5] (_5120),
        .\y[6] (_5121),
        .\y[7] (_5122),
        .\y[8] (_5123),
        .\y[9] (_5124),
        .\y[10] (_5125),
        .\y[11] (_5126),
        .\y[12] (_5127),
        .\y[13] (_5128),
        .\y[14] (_5129),
        .\y[15] (_5130)
    );
    swap u75 (
        .\a[0] (_4985),
        .\a[1] (_4986),
        .\a[2] (_4987),
        .\a[3] (_4988),
        .\a[4] (_4989),
        .\a[5] (_4990),
        .\a[6] (_4991),
        .\a[7] (_4992),
        .\a[8] (_4993),
        .\a[9] (_4994),
        .\a[10] (_4995),
        .\a[11] (_4996),
        .\a[12] (_4997),
        .\a[13] (_4998),
        .\a[14] (_4999),
        .\a[15] (_5000),
        .\b[0] (_5050),
        .\b[1] (_5051),
        .\b[2] (_5052),
        .\b[3] (_5053),
        .\b[4] (_5054),
        .\b[5] (_5055),
        .\b[6] (_5056),
        .\b[7] (_5057),
        .\b[8] (_5058),
        .\b[9] (_5059),
        .\b[10] (_5060),
        .\b[11] (_5061),
        .\b[12] (_5062),
        .\b[13] (_5063),
        .\b[14] (_5064),
        .\b[15] (_5065),
        .\x[0] (_5164),
        .\x[1] (_5165),
        .\x[2] (_5166),
        .\x[3] (_5167),
        .\x[4] (_5168),
        .\x[5] (_5169),
        .\x[6] (_5170),
        .\x[7] (_5171),
        .\x[8] (_5172),
        .\x[9] (_5173),
        .\x[10] (_5174),
        .\x[11] (_5175),
        .\x[12] (_5176),
        .\x[13] (_5177),
        .\x[14] (_5178),
        .\x[15] (_5179),
        .\y[0] (_5180),
        .\y[1] (_5181),
        .\y[2] (_5182),
        .\y[3] (_5183),
        .\y[4] (_5184),
        .\y[5] (_5185),
        .\y[6] (_5186),
        .\y[7] (_5187),
        .\y[8] (_5188),
        .\y[9] (_5189),
        .\y[10] (_5190),
        .\y[11] (_5191),
        .\y[12] (_5192),
        .\y[13] (_5193),
        .\y[14] (_5194),
        .\y[15] (_5195)
    );
    swap u76 (
        .\a[0] (_4725),
        .\a[1] (_4726),
        .\a[2] (_4727),
        .\a[3] (_4728),
        .\a[4] (_4729),
        .\a[5] (_4730),
        .\a[6] (_4731),
        .\a[7] (_4732),
        .\a[8] (_4733),
        .\a[9] (_4734),
        .\a[10] (_4735),
        .\a[11] (_4736),
        .\a[12] (_4737),
        .\a[13] (_4738),
        .\a[14] (_4739),
        .\a[15] (_4740),
        .\b[0] (_4855),
        .\b[1] (_4856),
        .\b[2] (_4857),
        .\b[3] (_4858),
        .\b[4] (_4859),
        .\b[5] (_4860),
        .\b[6] (_4861),
        .\b[7] (_4862),
        .\b[8] (_4863),
        .\b[9] (_4864),
        .\b[10] (_4865),
        .\b[11] (_4866),
        .\b[12] (_4867),
        .\b[13] (_4868),
        .\b[14] (_4869),
        .\b[15] (_4870),
        .\x[0] (_5229),
        .\x[1] (_5230),
        .\x[2] (_5231),
        .\x[3] (_5232),
        .\x[4] (_5233),
        .\x[5] (_5234),
        .\x[6] (_5235),
        .\x[7] (_5236),
        .\x[8] (_5237),
        .\x[9] (_5238),
        .\x[10] (_5239),
        .\x[11] (_5240),
        .\x[12] (_5241),
        .\x[13] (_5242),
        .\x[14] (_5243),
        .\x[15] (_5244),
        .\y[0] (_5245),
        .\y[1] (_5246),
        .\y[2] (_5247),
        .\y[3] (_5248),
        .\y[4] (_5249),
        .\y[5] (_5250),
        .\y[6] (_5251),
        .\y[7] (_5252),
        .\y[8] (_5253),
        .\y[9] (_5254),
        .\y[10] (_5255),
        .\y[11] (_5256),
        .\y[12] (_5257),
        .\y[13] (_5258),
        .\y[14] (_5259),
        .\y[15] (_5260)
    );
    swap u77 (
        .\a[0] (_4790),
        .\a[1] (_4791),
        .\a[2] (_4792),
        .\a[3] (_4793),
        .\a[4] (_4794),
        .\a[5] (_4795),
        .\a[6] (_4796),
        .\a[7] (_4797),
        .\a[8] (_4798),
        .\a[9] (_4799),
        .\a[10] (_4800),
        .\a[11] (_4801),
        .\a[12] (_4802),
        .\a[13] (_4803),
        .\a[14] (_4804),
        .\a[15] (_4805),
        .\b[0] (_4920),
        .\b[1] (_4921),
        .\b[2] (_4922),
        .\b[3] (_4923),
        .\b[4] (_4924),
        .\b[5] (_4925),
        .\b[6] (_4926),
        .\b[7] (_4927),
        .\b[8] (_4928),
        .\b[9] (_4929),
        .\b[10] (_4930),
        .\b[11] (_4931),
        .\b[12] (_4932),
        .\b[13] (_4933),
        .\b[14] (_4934),
        .\b[15] (_4935),
        .\x[0] (_5294),
        .\x[1] (_5295),
        .\x[2] (_5296),
        .\x[3] (_5297),
        .\x[4] (_5298),
        .\x[5] (_5299),
        .\x[6] (_5300),
        .\x[7] (_5301),
        .\x[8] (_5302),
        .\x[9] (_5303),
        .\x[10] (_5304),
        .\x[11] (_5305),
        .\x[12] (_5306),
        .\x[13] (_5307),
        .\x[14] (_5308),
        .\x[15] (_5309),
        .\y[0] (_5310),
        .\y[1] (_5311),
        .\y[2] (_5312),
        .\y[3] (_5313),
        .\y[4] (_5314),
        .\y[5] (_5315),
        .\y[6] (_5316),
        .\y[7] (_5317),
        .\y[8] (_5318),
        .\y[9] (_5319),
        .\y[10] (_5320),
        .\y[11] (_5321),
        .\y[12] (_5322),
        .\y[13] (_5323),
        .\y[14] (_5324),
        .\y[15] (_5325)
    );
    swap u78 (
        .\a[0] (_5229),
        .\a[1] (_5230),
        .\a[2] (_5231),
        .\a[3] (_5232),
        .\a[4] (_5233),
        .\a[5] (_5234),
        .\a[6] (_5235),
        .\a[7] (_5236),
        .\a[8] (_5237),
        .\a[9] (_5238),
        .\a[10] (_5239),
        .\a[11] (_5240),
        .\a[12] (_5241),
        .\a[13] (_5242),
        .\a[14] (_5243),
        .\a[15] (_5244),
        .\b[0] (_5294),
        .\b[1] (_5295),
        .\b[2] (_5296),
        .\b[3] (_5297),
        .\b[4] (_5298),
        .\b[5] (_5299),
        .\b[6] (_5300),
        .\b[7] (_5301),
        .\b[8] (_5302),
        .\b[9] (_5303),
        .\b[10] (_5304),
        .\b[11] (_5305),
        .\b[12] (_5306),
        .\b[13] (_5307),
        .\b[14] (_5308),
        .\b[15] (_5309),
        .\x[0] (_5359),
        .\x[1] (_5360),
        .\x[2] (_5361),
        .\x[3] (_5362),
        .\x[4] (_5363),
        .\x[5] (_5364),
        .\x[6] (_5365),
        .\x[7] (_5366),
        .\x[8] (_5367),
        .\x[9] (_5368),
        .\x[10] (_5369),
        .\x[11] (_5370),
        .\x[12] (_5371),
        .\x[13] (_5372),
        .\x[14] (_5373),
        .\x[15] (_5374),
        .\y[0] (_5375),
        .\y[1] (_5376),
        .\y[2] (_5377),
        .\y[3] (_5378),
        .\y[4] (_5379),
        .\y[5] (_5380),
        .\y[6] (_5381),
        .\y[7] (_5382),
        .\y[8] (_5383),
        .\y[9] (_5384),
        .\y[10] (_5385),
        .\y[11] (_5386),
        .\y[12] (_5387),
        .\y[13] (_5388),
        .\y[14] (_5389),
        .\y[15] (_5390)
    );
    swap u79 (
        .\a[0] (_5245),
        .\a[1] (_5246),
        .\a[2] (_5247),
        .\a[3] (_5248),
        .\a[4] (_5249),
        .\a[5] (_5250),
        .\a[6] (_5251),
        .\a[7] (_5252),
        .\a[8] (_5253),
        .\a[9] (_5254),
        .\a[10] (_5255),
        .\a[11] (_5256),
        .\a[12] (_5257),
        .\a[13] (_5258),
        .\a[14] (_5259),
        .\a[15] (_5260),
        .\b[0] (_5310),
        .\b[1] (_5311),
        .\b[2] (_5312),
        .\b[3] (_5313),
        .\b[4] (_5314),
        .\b[5] (_5315),
        .\b[6] (_5316),
        .\b[7] (_5317),
        .\b[8] (_5318),
        .\b[9] (_5319),
        .\b[10] (_5320),
        .\b[11] (_5321),
        .\b[12] (_5322),
        .\b[13] (_5323),
        .\b[14] (_5324),
        .\b[15] (_5325),
        .\x[0] (_5424),
        .\x[1] (_5425),
        .\x[2] (_5426),
        .\x[3] (_5427),
        .\x[4] (_5428),
        .\x[5] (_5429),
        .\x[6] (_5430),
        .\x[7] (_5431),
        .\x[8] (_5432),
        .\x[9] (_5433),
        .\x[10] (_5434),
        .\x[11] (_5435),
        .\x[12] (_5436),
        .\x[13] (_5437),
        .\x[14] (_5438),
        .\x[15] (_5439),
        .\y[0] (_5440),
        .\y[1] (_5441),
        .\y[2] (_5442),
        .\y[3] (_5443),
        .\y[4] (_5444),
        .\y[5] (_5445),
        .\y[6] (_5446),
        .\y[7] (_5447),
        .\y[8] (_5448),
        .\y[9] (_5449),
        .\y[10] (_5450),
        .\y[11] (_5451),
        .\y[12] (_5452),
        .\y[13] (_5453),
        .\y[14] (_5454),
        .\y[15] (_5455)
    );
    always @(posedge clk) begin
        \a_sorted[0][0]  <= \a_sorted[0][0]_ns ;
        \a_sorted[0][1]  <= \a_sorted[0][1]_ns ;
        \a_sorted[0][2]  <= \a_sorted[0][2]_ns ;
        \a_sorted[0][3]  <= \a_sorted[0][3]_ns ;
        \a_sorted[0][4]  <= \a_sorted[0][4]_ns ;
        \a_sorted[0][5]  <= \a_sorted[0][5]_ns ;
        \a_sorted[0][6]  <= \a_sorted[0][6]_ns ;
        \a_sorted[0][7]  <= \a_sorted[0][7]_ns ;
        \a_sorted[0][8]  <= \a_sorted[0][8]_ns ;
        \a_sorted[0][9]  <= \a_sorted[0][9]_ns ;
        \a_sorted[0][10]  <= \a_sorted[0][10]_ns ;
        \a_sorted[0][11]  <= \a_sorted[0][11]_ns ;
        \a_sorted[0][12]  <= \a_sorted[0][12]_ns ;
        \a_sorted[0][13]  <= \a_sorted[0][13]_ns ;
        \a_sorted[0][14]  <= \a_sorted[0][14]_ns ;
        \a_sorted[0][15]  <= \a_sorted[0][15]_ns ;
        \a_sorted[1][0]  <= \a_sorted[1][0]_ns ;
        \a_sorted[1][1]  <= \a_sorted[1][1]_ns ;
        \a_sorted[1][2]  <= \a_sorted[1][2]_ns ;
        \a_sorted[1][3]  <= \a_sorted[1][3]_ns ;
        \a_sorted[1][4]  <= \a_sorted[1][4]_ns ;
        \a_sorted[1][5]  <= \a_sorted[1][5]_ns ;
        \a_sorted[1][6]  <= \a_sorted[1][6]_ns ;
        \a_sorted[1][7]  <= \a_sorted[1][7]_ns ;
        \a_sorted[1][8]  <= \a_sorted[1][8]_ns ;
        \a_sorted[1][9]  <= \a_sorted[1][9]_ns ;
        \a_sorted[1][10]  <= \a_sorted[1][10]_ns ;
        \a_sorted[1][11]  <= \a_sorted[1][11]_ns ;
        \a_sorted[1][12]  <= \a_sorted[1][12]_ns ;
        \a_sorted[1][13]  <= \a_sorted[1][13]_ns ;
        \a_sorted[1][14]  <= \a_sorted[1][14]_ns ;
        \a_sorted[1][15]  <= \a_sorted[1][15]_ns ;
        \a_sorted[2][0]  <= \a_sorted[2][0]_ns ;
        \a_sorted[2][1]  <= \a_sorted[2][1]_ns ;
        \a_sorted[2][2]  <= \a_sorted[2][2]_ns ;
        \a_sorted[2][3]  <= \a_sorted[2][3]_ns ;
        \a_sorted[2][4]  <= \a_sorted[2][4]_ns ;
        \a_sorted[2][5]  <= \a_sorted[2][5]_ns ;
        \a_sorted[2][6]  <= \a_sorted[2][6]_ns ;
        \a_sorted[2][7]  <= \a_sorted[2][7]_ns ;
        \a_sorted[2][8]  <= \a_sorted[2][8]_ns ;
        \a_sorted[2][9]  <= \a_sorted[2][9]_ns ;
        \a_sorted[2][10]  <= \a_sorted[2][10]_ns ;
        \a_sorted[2][11]  <= \a_sorted[2][11]_ns ;
        \a_sorted[2][12]  <= \a_sorted[2][12]_ns ;
        \a_sorted[2][13]  <= \a_sorted[2][13]_ns ;
        \a_sorted[2][14]  <= \a_sorted[2][14]_ns ;
        \a_sorted[2][15]  <= \a_sorted[2][15]_ns ;
        \a_sorted[3][0]  <= \a_sorted[3][0]_ns ;
        \a_sorted[3][1]  <= \a_sorted[3][1]_ns ;
        \a_sorted[3][2]  <= \a_sorted[3][2]_ns ;
        \a_sorted[3][3]  <= \a_sorted[3][3]_ns ;
        \a_sorted[3][4]  <= \a_sorted[3][4]_ns ;
        \a_sorted[3][5]  <= \a_sorted[3][5]_ns ;
        \a_sorted[3][6]  <= \a_sorted[3][6]_ns ;
        \a_sorted[3][7]  <= \a_sorted[3][7]_ns ;
        \a_sorted[3][8]  <= \a_sorted[3][8]_ns ;
        \a_sorted[3][9]  <= \a_sorted[3][9]_ns ;
        \a_sorted[3][10]  <= \a_sorted[3][10]_ns ;
        \a_sorted[3][11]  <= \a_sorted[3][11]_ns ;
        \a_sorted[3][12]  <= \a_sorted[3][12]_ns ;
        \a_sorted[3][13]  <= \a_sorted[3][13]_ns ;
        \a_sorted[3][14]  <= \a_sorted[3][14]_ns ;
        \a_sorted[3][15]  <= \a_sorted[3][15]_ns ;
        \a_sorted[4][0]  <= \a_sorted[4][0]_ns ;
        \a_sorted[4][1]  <= \a_sorted[4][1]_ns ;
        \a_sorted[4][2]  <= \a_sorted[4][2]_ns ;
        \a_sorted[4][3]  <= \a_sorted[4][3]_ns ;
        \a_sorted[4][4]  <= \a_sorted[4][4]_ns ;
        \a_sorted[4][5]  <= \a_sorted[4][5]_ns ;
        \a_sorted[4][6]  <= \a_sorted[4][6]_ns ;
        \a_sorted[4][7]  <= \a_sorted[4][7]_ns ;
        \a_sorted[4][8]  <= \a_sorted[4][8]_ns ;
        \a_sorted[4][9]  <= \a_sorted[4][9]_ns ;
        \a_sorted[4][10]  <= \a_sorted[4][10]_ns ;
        \a_sorted[4][11]  <= \a_sorted[4][11]_ns ;
        \a_sorted[4][12]  <= \a_sorted[4][12]_ns ;
        \a_sorted[4][13]  <= \a_sorted[4][13]_ns ;
        \a_sorted[4][14]  <= \a_sorted[4][14]_ns ;
        \a_sorted[4][15]  <= \a_sorted[4][15]_ns ;
        \a_sorted[5][0]  <= \a_sorted[5][0]_ns ;
        \a_sorted[5][1]  <= \a_sorted[5][1]_ns ;
        \a_sorted[5][2]  <= \a_sorted[5][2]_ns ;
        \a_sorted[5][3]  <= \a_sorted[5][3]_ns ;
        \a_sorted[5][4]  <= \a_sorted[5][4]_ns ;
        \a_sorted[5][5]  <= \a_sorted[5][5]_ns ;
        \a_sorted[5][6]  <= \a_sorted[5][6]_ns ;
        \a_sorted[5][7]  <= \a_sorted[5][7]_ns ;
        \a_sorted[5][8]  <= \a_sorted[5][8]_ns ;
        \a_sorted[5][9]  <= \a_sorted[5][9]_ns ;
        \a_sorted[5][10]  <= \a_sorted[5][10]_ns ;
        \a_sorted[5][11]  <= \a_sorted[5][11]_ns ;
        \a_sorted[5][12]  <= \a_sorted[5][12]_ns ;
        \a_sorted[5][13]  <= \a_sorted[5][13]_ns ;
        \a_sorted[5][14]  <= \a_sorted[5][14]_ns ;
        \a_sorted[5][15]  <= \a_sorted[5][15]_ns ;
        \a_sorted[6][0]  <= \a_sorted[6][0]_ns ;
        \a_sorted[6][1]  <= \a_sorted[6][1]_ns ;
        \a_sorted[6][2]  <= \a_sorted[6][2]_ns ;
        \a_sorted[6][3]  <= \a_sorted[6][3]_ns ;
        \a_sorted[6][4]  <= \a_sorted[6][4]_ns ;
        \a_sorted[6][5]  <= \a_sorted[6][5]_ns ;
        \a_sorted[6][6]  <= \a_sorted[6][6]_ns ;
        \a_sorted[6][7]  <= \a_sorted[6][7]_ns ;
        \a_sorted[6][8]  <= \a_sorted[6][8]_ns ;
        \a_sorted[6][9]  <= \a_sorted[6][9]_ns ;
        \a_sorted[6][10]  <= \a_sorted[6][10]_ns ;
        \a_sorted[6][11]  <= \a_sorted[6][11]_ns ;
        \a_sorted[6][12]  <= \a_sorted[6][12]_ns ;
        \a_sorted[6][13]  <= \a_sorted[6][13]_ns ;
        \a_sorted[6][14]  <= \a_sorted[6][14]_ns ;
        \a_sorted[6][15]  <= \a_sorted[6][15]_ns ;
        \a_sorted[7][0]  <= \a_sorted[7][0]_ns ;
        \a_sorted[7][1]  <= \a_sorted[7][1]_ns ;
        \a_sorted[7][2]  <= \a_sorted[7][2]_ns ;
        \a_sorted[7][3]  <= \a_sorted[7][3]_ns ;
        \a_sorted[7][4]  <= \a_sorted[7][4]_ns ;
        \a_sorted[7][5]  <= \a_sorted[7][5]_ns ;
        \a_sorted[7][6]  <= \a_sorted[7][6]_ns ;
        \a_sorted[7][7]  <= \a_sorted[7][7]_ns ;
        \a_sorted[7][8]  <= \a_sorted[7][8]_ns ;
        \a_sorted[7][9]  <= \a_sorted[7][9]_ns ;
        \a_sorted[7][10]  <= \a_sorted[7][10]_ns ;
        \a_sorted[7][11]  <= \a_sorted[7][11]_ns ;
        \a_sorted[7][12]  <= \a_sorted[7][12]_ns ;
        \a_sorted[7][13]  <= \a_sorted[7][13]_ns ;
        \a_sorted[7][14]  <= \a_sorted[7][14]_ns ;
        \a_sorted[7][15]  <= \a_sorted[7][15]_ns ;
        \a_sorted[8][0]  <= \a_sorted[8][0]_ns ;
        \a_sorted[8][1]  <= \a_sorted[8][1]_ns ;
        \a_sorted[8][2]  <= \a_sorted[8][2]_ns ;
        \a_sorted[8][3]  <= \a_sorted[8][3]_ns ;
        \a_sorted[8][4]  <= \a_sorted[8][4]_ns ;
        \a_sorted[8][5]  <= \a_sorted[8][5]_ns ;
        \a_sorted[8][6]  <= \a_sorted[8][6]_ns ;
        \a_sorted[8][7]  <= \a_sorted[8][7]_ns ;
        \a_sorted[8][8]  <= \a_sorted[8][8]_ns ;
        \a_sorted[8][9]  <= \a_sorted[8][9]_ns ;
        \a_sorted[8][10]  <= \a_sorted[8][10]_ns ;
        \a_sorted[8][11]  <= \a_sorted[8][11]_ns ;
        \a_sorted[8][12]  <= \a_sorted[8][12]_ns ;
        \a_sorted[8][13]  <= \a_sorted[8][13]_ns ;
        \a_sorted[8][14]  <= \a_sorted[8][14]_ns ;
        \a_sorted[8][15]  <= \a_sorted[8][15]_ns ;
        \a_sorted[9][0]  <= \a_sorted[9][0]_ns ;
        \a_sorted[9][1]  <= \a_sorted[9][1]_ns ;
        \a_sorted[9][2]  <= \a_sorted[9][2]_ns ;
        \a_sorted[9][3]  <= \a_sorted[9][3]_ns ;
        \a_sorted[9][4]  <= \a_sorted[9][4]_ns ;
        \a_sorted[9][5]  <= \a_sorted[9][5]_ns ;
        \a_sorted[9][6]  <= \a_sorted[9][6]_ns ;
        \a_sorted[9][7]  <= \a_sorted[9][7]_ns ;
        \a_sorted[9][8]  <= \a_sorted[9][8]_ns ;
        \a_sorted[9][9]  <= \a_sorted[9][9]_ns ;
        \a_sorted[9][10]  <= \a_sorted[9][10]_ns ;
        \a_sorted[9][11]  <= \a_sorted[9][11]_ns ;
        \a_sorted[9][12]  <= \a_sorted[9][12]_ns ;
        \a_sorted[9][13]  <= \a_sorted[9][13]_ns ;
        \a_sorted[9][14]  <= \a_sorted[9][14]_ns ;
        \a_sorted[9][15]  <= \a_sorted[9][15]_ns ;
        \a_sorted[10][0]  <= \a_sorted[10][0]_ns ;
        \a_sorted[10][1]  <= \a_sorted[10][1]_ns ;
        \a_sorted[10][2]  <= \a_sorted[10][2]_ns ;
        \a_sorted[10][3]  <= \a_sorted[10][3]_ns ;
        \a_sorted[10][4]  <= \a_sorted[10][4]_ns ;
        \a_sorted[10][5]  <= \a_sorted[10][5]_ns ;
        \a_sorted[10][6]  <= \a_sorted[10][6]_ns ;
        \a_sorted[10][7]  <= \a_sorted[10][7]_ns ;
        \a_sorted[10][8]  <= \a_sorted[10][8]_ns ;
        \a_sorted[10][9]  <= \a_sorted[10][9]_ns ;
        \a_sorted[10][10]  <= \a_sorted[10][10]_ns ;
        \a_sorted[10][11]  <= \a_sorted[10][11]_ns ;
        \a_sorted[10][12]  <= \a_sorted[10][12]_ns ;
        \a_sorted[10][13]  <= \a_sorted[10][13]_ns ;
        \a_sorted[10][14]  <= \a_sorted[10][14]_ns ;
        \a_sorted[10][15]  <= \a_sorted[10][15]_ns ;
        \a_sorted[11][0]  <= \a_sorted[11][0]_ns ;
        \a_sorted[11][1]  <= \a_sorted[11][1]_ns ;
        \a_sorted[11][2]  <= \a_sorted[11][2]_ns ;
        \a_sorted[11][3]  <= \a_sorted[11][3]_ns ;
        \a_sorted[11][4]  <= \a_sorted[11][4]_ns ;
        \a_sorted[11][5]  <= \a_sorted[11][5]_ns ;
        \a_sorted[11][6]  <= \a_sorted[11][6]_ns ;
        \a_sorted[11][7]  <= \a_sorted[11][7]_ns ;
        \a_sorted[11][8]  <= \a_sorted[11][8]_ns ;
        \a_sorted[11][9]  <= \a_sorted[11][9]_ns ;
        \a_sorted[11][10]  <= \a_sorted[11][10]_ns ;
        \a_sorted[11][11]  <= \a_sorted[11][11]_ns ;
        \a_sorted[11][12]  <= \a_sorted[11][12]_ns ;
        \a_sorted[11][13]  <= \a_sorted[11][13]_ns ;
        \a_sorted[11][14]  <= \a_sorted[11][14]_ns ;
        \a_sorted[11][15]  <= \a_sorted[11][15]_ns ;
        \a_sorted[12][0]  <= \a_sorted[12][0]_ns ;
        \a_sorted[12][1]  <= \a_sorted[12][1]_ns ;
        \a_sorted[12][2]  <= \a_sorted[12][2]_ns ;
        \a_sorted[12][3]  <= \a_sorted[12][3]_ns ;
        \a_sorted[12][4]  <= \a_sorted[12][4]_ns ;
        \a_sorted[12][5]  <= \a_sorted[12][5]_ns ;
        \a_sorted[12][6]  <= \a_sorted[12][6]_ns ;
        \a_sorted[12][7]  <= \a_sorted[12][7]_ns ;
        \a_sorted[12][8]  <= \a_sorted[12][8]_ns ;
        \a_sorted[12][9]  <= \a_sorted[12][9]_ns ;
        \a_sorted[12][10]  <= \a_sorted[12][10]_ns ;
        \a_sorted[12][11]  <= \a_sorted[12][11]_ns ;
        \a_sorted[12][12]  <= \a_sorted[12][12]_ns ;
        \a_sorted[12][13]  <= \a_sorted[12][13]_ns ;
        \a_sorted[12][14]  <= \a_sorted[12][14]_ns ;
        \a_sorted[12][15]  <= \a_sorted[12][15]_ns ;
        \a_sorted[13][0]  <= \a_sorted[13][0]_ns ;
        \a_sorted[13][1]  <= \a_sorted[13][1]_ns ;
        \a_sorted[13][2]  <= \a_sorted[13][2]_ns ;
        \a_sorted[13][3]  <= \a_sorted[13][3]_ns ;
        \a_sorted[13][4]  <= \a_sorted[13][4]_ns ;
        \a_sorted[13][5]  <= \a_sorted[13][5]_ns ;
        \a_sorted[13][6]  <= \a_sorted[13][6]_ns ;
        \a_sorted[13][7]  <= \a_sorted[13][7]_ns ;
        \a_sorted[13][8]  <= \a_sorted[13][8]_ns ;
        \a_sorted[13][9]  <= \a_sorted[13][9]_ns ;
        \a_sorted[13][10]  <= \a_sorted[13][10]_ns ;
        \a_sorted[13][11]  <= \a_sorted[13][11]_ns ;
        \a_sorted[13][12]  <= \a_sorted[13][12]_ns ;
        \a_sorted[13][13]  <= \a_sorted[13][13]_ns ;
        \a_sorted[13][14]  <= \a_sorted[13][14]_ns ;
        \a_sorted[13][15]  <= \a_sorted[13][15]_ns ;
        \a_sorted[14][0]  <= \a_sorted[14][0]_ns ;
        \a_sorted[14][1]  <= \a_sorted[14][1]_ns ;
        \a_sorted[14][2]  <= \a_sorted[14][2]_ns ;
        \a_sorted[14][3]  <= \a_sorted[14][3]_ns ;
        \a_sorted[14][4]  <= \a_sorted[14][4]_ns ;
        \a_sorted[14][5]  <= \a_sorted[14][5]_ns ;
        \a_sorted[14][6]  <= \a_sorted[14][6]_ns ;
        \a_sorted[14][7]  <= \a_sorted[14][7]_ns ;
        \a_sorted[14][8]  <= \a_sorted[14][8]_ns ;
        \a_sorted[14][9]  <= \a_sorted[14][9]_ns ;
        \a_sorted[14][10]  <= \a_sorted[14][10]_ns ;
        \a_sorted[14][11]  <= \a_sorted[14][11]_ns ;
        \a_sorted[14][12]  <= \a_sorted[14][12]_ns ;
        \a_sorted[14][13]  <= \a_sorted[14][13]_ns ;
        \a_sorted[14][14]  <= \a_sorted[14][14]_ns ;
        \a_sorted[14][15]  <= \a_sorted[14][15]_ns ;
        \a_sorted[15][0]  <= \a_sorted[15][0]_ns ;
        \a_sorted[15][1]  <= \a_sorted[15][1]_ns ;
        \a_sorted[15][2]  <= \a_sorted[15][2]_ns ;
        \a_sorted[15][3]  <= \a_sorted[15][3]_ns ;
        \a_sorted[15][4]  <= \a_sorted[15][4]_ns ;
        \a_sorted[15][5]  <= \a_sorted[15][5]_ns ;
        \a_sorted[15][6]  <= \a_sorted[15][6]_ns ;
        \a_sorted[15][7]  <= \a_sorted[15][7]_ns ;
        \a_sorted[15][8]  <= \a_sorted[15][8]_ns ;
        \a_sorted[15][9]  <= \a_sorted[15][9]_ns ;
        \a_sorted[15][10]  <= \a_sorted[15][10]_ns ;
        \a_sorted[15][11]  <= \a_sorted[15][11]_ns ;
        \a_sorted[15][12]  <= \a_sorted[15][12]_ns ;
        \a_sorted[15][13]  <= \a_sorted[15][13]_ns ;
        \a_sorted[15][14]  <= \a_sorted[15][14]_ns ;
        \a_sorted[15][15]  <= \a_sorted[15][15]_ns ;
    end
endmodule

